module ProcessorTopLevel(
  input   clock,
  input   reset
);
endmodule
