module InstrMemoryTest(
  input         clock,
  input         reset,
  input  [9:0]  io_addr,
  output [31:0] io_dataOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] dataReg; // @[InstrMemoryTest.scala 20:24]
  wire [31:0] _GEN_8 = 10'h8 == io_addr ? 32'h0 : 32'h13; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_9 = 10'h9 == io_addr ? 32'h0 : _GEN_8; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_10 = 10'ha == io_addr ? 32'h0 : _GEN_9; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_11 = 10'hb == io_addr ? 32'h0 : _GEN_10; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_12 = 10'hc == io_addr ? 32'h0 : _GEN_11; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_13 = 10'hd == io_addr ? 32'h0 : _GEN_12; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_14 = 10'he == io_addr ? 32'h0 : _GEN_13; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_15 = 10'hf == io_addr ? 32'h0 : _GEN_14; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_16 = 10'h10 == io_addr ? 32'h0 : _GEN_15; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_17 = 10'h11 == io_addr ? 32'h0 : _GEN_16; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_18 = 10'h12 == io_addr ? 32'h0 : _GEN_17; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_19 = 10'h13 == io_addr ? 32'h0 : _GEN_18; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_20 = 10'h14 == io_addr ? 32'h0 : _GEN_19; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_21 = 10'h15 == io_addr ? 32'h0 : _GEN_20; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_22 = 10'h16 == io_addr ? 32'h0 : _GEN_21; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_23 = 10'h17 == io_addr ? 32'h0 : _GEN_22; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_24 = 10'h18 == io_addr ? 32'h0 : _GEN_23; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_25 = 10'h19 == io_addr ? 32'h0 : _GEN_24; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_26 = 10'h1a == io_addr ? 32'h0 : _GEN_25; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_27 = 10'h1b == io_addr ? 32'h0 : _GEN_26; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_28 = 10'h1c == io_addr ? 32'h0 : _GEN_27; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_29 = 10'h1d == io_addr ? 32'h0 : _GEN_28; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_30 = 10'h1e == io_addr ? 32'h0 : _GEN_29; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_31 = 10'h1f == io_addr ? 32'h0 : _GEN_30; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_32 = 10'h20 == io_addr ? 32'h0 : _GEN_31; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_33 = 10'h21 == io_addr ? 32'h0 : _GEN_32; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_34 = 10'h22 == io_addr ? 32'h0 : _GEN_33; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_35 = 10'h23 == io_addr ? 32'h0 : _GEN_34; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_36 = 10'h24 == io_addr ? 32'h0 : _GEN_35; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_37 = 10'h25 == io_addr ? 32'h0 : _GEN_36; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_38 = 10'h26 == io_addr ? 32'h0 : _GEN_37; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_39 = 10'h27 == io_addr ? 32'h0 : _GEN_38; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_40 = 10'h28 == io_addr ? 32'h0 : _GEN_39; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_41 = 10'h29 == io_addr ? 32'h0 : _GEN_40; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_42 = 10'h2a == io_addr ? 32'h0 : _GEN_41; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_43 = 10'h2b == io_addr ? 32'h0 : _GEN_42; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_44 = 10'h2c == io_addr ? 32'h0 : _GEN_43; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_45 = 10'h2d == io_addr ? 32'h0 : _GEN_44; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_46 = 10'h2e == io_addr ? 32'h0 : _GEN_45; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_47 = 10'h2f == io_addr ? 32'h0 : _GEN_46; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_48 = 10'h30 == io_addr ? 32'h0 : _GEN_47; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_49 = 10'h31 == io_addr ? 32'h0 : _GEN_48; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_50 = 10'h32 == io_addr ? 32'h0 : _GEN_49; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_51 = 10'h33 == io_addr ? 32'h0 : _GEN_50; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_52 = 10'h34 == io_addr ? 32'h0 : _GEN_51; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_53 = 10'h35 == io_addr ? 32'h0 : _GEN_52; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_54 = 10'h36 == io_addr ? 32'h0 : _GEN_53; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_55 = 10'h37 == io_addr ? 32'h0 : _GEN_54; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_56 = 10'h38 == io_addr ? 32'h0 : _GEN_55; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_57 = 10'h39 == io_addr ? 32'h0 : _GEN_56; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_58 = 10'h3a == io_addr ? 32'h0 : _GEN_57; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_59 = 10'h3b == io_addr ? 32'h0 : _GEN_58; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_60 = 10'h3c == io_addr ? 32'h0 : _GEN_59; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_61 = 10'h3d == io_addr ? 32'h0 : _GEN_60; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_62 = 10'h3e == io_addr ? 32'h0 : _GEN_61; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_63 = 10'h3f == io_addr ? 32'h0 : _GEN_62; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_64 = 10'h40 == io_addr ? 32'h0 : _GEN_63; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_65 = 10'h41 == io_addr ? 32'h0 : _GEN_64; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_66 = 10'h42 == io_addr ? 32'h0 : _GEN_65; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_67 = 10'h43 == io_addr ? 32'h0 : _GEN_66; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_68 = 10'h44 == io_addr ? 32'h0 : _GEN_67; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_69 = 10'h45 == io_addr ? 32'h0 : _GEN_68; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_70 = 10'h46 == io_addr ? 32'h0 : _GEN_69; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_71 = 10'h47 == io_addr ? 32'h0 : _GEN_70; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_72 = 10'h48 == io_addr ? 32'h0 : _GEN_71; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_73 = 10'h49 == io_addr ? 32'h0 : _GEN_72; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_74 = 10'h4a == io_addr ? 32'h0 : _GEN_73; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_75 = 10'h4b == io_addr ? 32'h0 : _GEN_74; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_76 = 10'h4c == io_addr ? 32'h0 : _GEN_75; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_77 = 10'h4d == io_addr ? 32'h0 : _GEN_76; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_78 = 10'h4e == io_addr ? 32'h0 : _GEN_77; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_79 = 10'h4f == io_addr ? 32'h0 : _GEN_78; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_80 = 10'h50 == io_addr ? 32'h0 : _GEN_79; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_81 = 10'h51 == io_addr ? 32'h0 : _GEN_80; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_82 = 10'h52 == io_addr ? 32'h0 : _GEN_81; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_83 = 10'h53 == io_addr ? 32'h0 : _GEN_82; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_84 = 10'h54 == io_addr ? 32'h0 : _GEN_83; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_85 = 10'h55 == io_addr ? 32'h0 : _GEN_84; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_86 = 10'h56 == io_addr ? 32'h0 : _GEN_85; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_87 = 10'h57 == io_addr ? 32'h0 : _GEN_86; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_88 = 10'h58 == io_addr ? 32'h0 : _GEN_87; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_89 = 10'h59 == io_addr ? 32'h0 : _GEN_88; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_90 = 10'h5a == io_addr ? 32'h0 : _GEN_89; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_91 = 10'h5b == io_addr ? 32'h0 : _GEN_90; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_92 = 10'h5c == io_addr ? 32'h0 : _GEN_91; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_93 = 10'h5d == io_addr ? 32'h0 : _GEN_92; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_94 = 10'h5e == io_addr ? 32'h0 : _GEN_93; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_95 = 10'h5f == io_addr ? 32'h0 : _GEN_94; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_96 = 10'h60 == io_addr ? 32'h0 : _GEN_95; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_97 = 10'h61 == io_addr ? 32'h0 : _GEN_96; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_98 = 10'h62 == io_addr ? 32'h0 : _GEN_97; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_99 = 10'h63 == io_addr ? 32'h0 : _GEN_98; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_100 = 10'h64 == io_addr ? 32'h0 : _GEN_99; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_101 = 10'h65 == io_addr ? 32'h0 : _GEN_100; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_102 = 10'h66 == io_addr ? 32'h0 : _GEN_101; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_103 = 10'h67 == io_addr ? 32'h0 : _GEN_102; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_104 = 10'h68 == io_addr ? 32'h0 : _GEN_103; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_105 = 10'h69 == io_addr ? 32'h0 : _GEN_104; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_106 = 10'h6a == io_addr ? 32'h0 : _GEN_105; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_107 = 10'h6b == io_addr ? 32'h0 : _GEN_106; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_108 = 10'h6c == io_addr ? 32'h0 : _GEN_107; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_109 = 10'h6d == io_addr ? 32'h0 : _GEN_108; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_110 = 10'h6e == io_addr ? 32'h0 : _GEN_109; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_111 = 10'h6f == io_addr ? 32'h0 : _GEN_110; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_112 = 10'h70 == io_addr ? 32'h0 : _GEN_111; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_113 = 10'h71 == io_addr ? 32'h0 : _GEN_112; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_114 = 10'h72 == io_addr ? 32'h0 : _GEN_113; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_115 = 10'h73 == io_addr ? 32'h0 : _GEN_114; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_116 = 10'h74 == io_addr ? 32'h0 : _GEN_115; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_117 = 10'h75 == io_addr ? 32'h0 : _GEN_116; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_118 = 10'h76 == io_addr ? 32'h0 : _GEN_117; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_119 = 10'h77 == io_addr ? 32'h0 : _GEN_118; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_120 = 10'h78 == io_addr ? 32'h0 : _GEN_119; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_121 = 10'h79 == io_addr ? 32'h0 : _GEN_120; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_122 = 10'h7a == io_addr ? 32'h0 : _GEN_121; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_123 = 10'h7b == io_addr ? 32'h0 : _GEN_122; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_124 = 10'h7c == io_addr ? 32'h0 : _GEN_123; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_125 = 10'h7d == io_addr ? 32'h0 : _GEN_124; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_126 = 10'h7e == io_addr ? 32'h0 : _GEN_125; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_127 = 10'h7f == io_addr ? 32'h0 : _GEN_126; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_128 = 10'h80 == io_addr ? 32'h0 : _GEN_127; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_129 = 10'h81 == io_addr ? 32'h0 : _GEN_128; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_130 = 10'h82 == io_addr ? 32'h0 : _GEN_129; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_131 = 10'h83 == io_addr ? 32'h0 : _GEN_130; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_132 = 10'h84 == io_addr ? 32'h0 : _GEN_131; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_133 = 10'h85 == io_addr ? 32'h0 : _GEN_132; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_134 = 10'h86 == io_addr ? 32'h0 : _GEN_133; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_135 = 10'h87 == io_addr ? 32'h0 : _GEN_134; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_136 = 10'h88 == io_addr ? 32'h0 : _GEN_135; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_137 = 10'h89 == io_addr ? 32'h0 : _GEN_136; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_138 = 10'h8a == io_addr ? 32'h0 : _GEN_137; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_139 = 10'h8b == io_addr ? 32'h0 : _GEN_138; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_140 = 10'h8c == io_addr ? 32'h0 : _GEN_139; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_141 = 10'h8d == io_addr ? 32'h0 : _GEN_140; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_142 = 10'h8e == io_addr ? 32'h0 : _GEN_141; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_143 = 10'h8f == io_addr ? 32'h0 : _GEN_142; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_144 = 10'h90 == io_addr ? 32'h0 : _GEN_143; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_145 = 10'h91 == io_addr ? 32'h0 : _GEN_144; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_146 = 10'h92 == io_addr ? 32'h0 : _GEN_145; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_147 = 10'h93 == io_addr ? 32'h0 : _GEN_146; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_148 = 10'h94 == io_addr ? 32'h0 : _GEN_147; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_149 = 10'h95 == io_addr ? 32'h0 : _GEN_148; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_150 = 10'h96 == io_addr ? 32'h0 : _GEN_149; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_151 = 10'h97 == io_addr ? 32'h0 : _GEN_150; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_152 = 10'h98 == io_addr ? 32'h0 : _GEN_151; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_153 = 10'h99 == io_addr ? 32'h0 : _GEN_152; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_154 = 10'h9a == io_addr ? 32'h0 : _GEN_153; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_155 = 10'h9b == io_addr ? 32'h0 : _GEN_154; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_156 = 10'h9c == io_addr ? 32'h0 : _GEN_155; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_157 = 10'h9d == io_addr ? 32'h0 : _GEN_156; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_158 = 10'h9e == io_addr ? 32'h0 : _GEN_157; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_159 = 10'h9f == io_addr ? 32'h0 : _GEN_158; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_160 = 10'ha0 == io_addr ? 32'h0 : _GEN_159; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_161 = 10'ha1 == io_addr ? 32'h0 : _GEN_160; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_162 = 10'ha2 == io_addr ? 32'h0 : _GEN_161; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_163 = 10'ha3 == io_addr ? 32'h0 : _GEN_162; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_164 = 10'ha4 == io_addr ? 32'h0 : _GEN_163; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_165 = 10'ha5 == io_addr ? 32'h0 : _GEN_164; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_166 = 10'ha6 == io_addr ? 32'h0 : _GEN_165; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_167 = 10'ha7 == io_addr ? 32'h0 : _GEN_166; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_168 = 10'ha8 == io_addr ? 32'h0 : _GEN_167; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_169 = 10'ha9 == io_addr ? 32'h0 : _GEN_168; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_170 = 10'haa == io_addr ? 32'h0 : _GEN_169; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_171 = 10'hab == io_addr ? 32'h0 : _GEN_170; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_172 = 10'hac == io_addr ? 32'h0 : _GEN_171; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_173 = 10'had == io_addr ? 32'h0 : _GEN_172; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_174 = 10'hae == io_addr ? 32'h0 : _GEN_173; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_175 = 10'haf == io_addr ? 32'h0 : _GEN_174; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_176 = 10'hb0 == io_addr ? 32'h0 : _GEN_175; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_177 = 10'hb1 == io_addr ? 32'h0 : _GEN_176; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_178 = 10'hb2 == io_addr ? 32'h0 : _GEN_177; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_179 = 10'hb3 == io_addr ? 32'h0 : _GEN_178; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_180 = 10'hb4 == io_addr ? 32'h0 : _GEN_179; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_181 = 10'hb5 == io_addr ? 32'h0 : _GEN_180; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_182 = 10'hb6 == io_addr ? 32'h0 : _GEN_181; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_183 = 10'hb7 == io_addr ? 32'h0 : _GEN_182; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_184 = 10'hb8 == io_addr ? 32'h0 : _GEN_183; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_185 = 10'hb9 == io_addr ? 32'h0 : _GEN_184; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_186 = 10'hba == io_addr ? 32'h0 : _GEN_185; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_187 = 10'hbb == io_addr ? 32'h0 : _GEN_186; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_188 = 10'hbc == io_addr ? 32'h0 : _GEN_187; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_189 = 10'hbd == io_addr ? 32'h0 : _GEN_188; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_190 = 10'hbe == io_addr ? 32'h0 : _GEN_189; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_191 = 10'hbf == io_addr ? 32'h0 : _GEN_190; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_192 = 10'hc0 == io_addr ? 32'h0 : _GEN_191; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_193 = 10'hc1 == io_addr ? 32'h0 : _GEN_192; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_194 = 10'hc2 == io_addr ? 32'h0 : _GEN_193; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_195 = 10'hc3 == io_addr ? 32'h0 : _GEN_194; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_196 = 10'hc4 == io_addr ? 32'h0 : _GEN_195; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_197 = 10'hc5 == io_addr ? 32'h0 : _GEN_196; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_198 = 10'hc6 == io_addr ? 32'h0 : _GEN_197; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_199 = 10'hc7 == io_addr ? 32'h0 : _GEN_198; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_200 = 10'hc8 == io_addr ? 32'h0 : _GEN_199; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_201 = 10'hc9 == io_addr ? 32'h0 : _GEN_200; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_202 = 10'hca == io_addr ? 32'h0 : _GEN_201; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_203 = 10'hcb == io_addr ? 32'h0 : _GEN_202; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_204 = 10'hcc == io_addr ? 32'h0 : _GEN_203; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_205 = 10'hcd == io_addr ? 32'h0 : _GEN_204; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_206 = 10'hce == io_addr ? 32'h0 : _GEN_205; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_207 = 10'hcf == io_addr ? 32'h0 : _GEN_206; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_208 = 10'hd0 == io_addr ? 32'h0 : _GEN_207; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_209 = 10'hd1 == io_addr ? 32'h0 : _GEN_208; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_210 = 10'hd2 == io_addr ? 32'h0 : _GEN_209; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_211 = 10'hd3 == io_addr ? 32'h0 : _GEN_210; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_212 = 10'hd4 == io_addr ? 32'h0 : _GEN_211; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_213 = 10'hd5 == io_addr ? 32'h0 : _GEN_212; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_214 = 10'hd6 == io_addr ? 32'h0 : _GEN_213; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_215 = 10'hd7 == io_addr ? 32'h0 : _GEN_214; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_216 = 10'hd8 == io_addr ? 32'h0 : _GEN_215; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_217 = 10'hd9 == io_addr ? 32'h0 : _GEN_216; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_218 = 10'hda == io_addr ? 32'h0 : _GEN_217; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_219 = 10'hdb == io_addr ? 32'h0 : _GEN_218; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_220 = 10'hdc == io_addr ? 32'h0 : _GEN_219; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_221 = 10'hdd == io_addr ? 32'h0 : _GEN_220; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_222 = 10'hde == io_addr ? 32'h0 : _GEN_221; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_223 = 10'hdf == io_addr ? 32'h0 : _GEN_222; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_224 = 10'he0 == io_addr ? 32'h0 : _GEN_223; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_225 = 10'he1 == io_addr ? 32'h0 : _GEN_224; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_226 = 10'he2 == io_addr ? 32'h0 : _GEN_225; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_227 = 10'he3 == io_addr ? 32'h0 : _GEN_226; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_228 = 10'he4 == io_addr ? 32'h0 : _GEN_227; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_229 = 10'he5 == io_addr ? 32'h0 : _GEN_228; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_230 = 10'he6 == io_addr ? 32'h0 : _GEN_229; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_231 = 10'he7 == io_addr ? 32'h0 : _GEN_230; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_232 = 10'he8 == io_addr ? 32'h0 : _GEN_231; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_233 = 10'he9 == io_addr ? 32'h0 : _GEN_232; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_234 = 10'hea == io_addr ? 32'h0 : _GEN_233; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_235 = 10'heb == io_addr ? 32'h0 : _GEN_234; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_236 = 10'hec == io_addr ? 32'h0 : _GEN_235; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_237 = 10'hed == io_addr ? 32'h0 : _GEN_236; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_238 = 10'hee == io_addr ? 32'h0 : _GEN_237; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_239 = 10'hef == io_addr ? 32'h0 : _GEN_238; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_240 = 10'hf0 == io_addr ? 32'h0 : _GEN_239; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_241 = 10'hf1 == io_addr ? 32'h0 : _GEN_240; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_242 = 10'hf2 == io_addr ? 32'h0 : _GEN_241; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_243 = 10'hf3 == io_addr ? 32'h0 : _GEN_242; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_244 = 10'hf4 == io_addr ? 32'h0 : _GEN_243; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_245 = 10'hf5 == io_addr ? 32'h0 : _GEN_244; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_246 = 10'hf6 == io_addr ? 32'h0 : _GEN_245; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_247 = 10'hf7 == io_addr ? 32'h0 : _GEN_246; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_248 = 10'hf8 == io_addr ? 32'h0 : _GEN_247; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_249 = 10'hf9 == io_addr ? 32'h0 : _GEN_248; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_250 = 10'hfa == io_addr ? 32'h0 : _GEN_249; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_251 = 10'hfb == io_addr ? 32'h0 : _GEN_250; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_252 = 10'hfc == io_addr ? 32'h0 : _GEN_251; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_253 = 10'hfd == io_addr ? 32'h0 : _GEN_252; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_254 = 10'hfe == io_addr ? 32'h0 : _GEN_253; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_255 = 10'hff == io_addr ? 32'h0 : _GEN_254; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_256 = 10'h100 == io_addr ? 32'h0 : _GEN_255; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_257 = 10'h101 == io_addr ? 32'h0 : _GEN_256; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_258 = 10'h102 == io_addr ? 32'h0 : _GEN_257; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_259 = 10'h103 == io_addr ? 32'h0 : _GEN_258; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_260 = 10'h104 == io_addr ? 32'h0 : _GEN_259; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_261 = 10'h105 == io_addr ? 32'h0 : _GEN_260; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_262 = 10'h106 == io_addr ? 32'h0 : _GEN_261; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_263 = 10'h107 == io_addr ? 32'h0 : _GEN_262; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_264 = 10'h108 == io_addr ? 32'h0 : _GEN_263; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_265 = 10'h109 == io_addr ? 32'h0 : _GEN_264; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_266 = 10'h10a == io_addr ? 32'h0 : _GEN_265; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_267 = 10'h10b == io_addr ? 32'h0 : _GEN_266; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_268 = 10'h10c == io_addr ? 32'h0 : _GEN_267; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_269 = 10'h10d == io_addr ? 32'h0 : _GEN_268; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_270 = 10'h10e == io_addr ? 32'h0 : _GEN_269; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_271 = 10'h10f == io_addr ? 32'h0 : _GEN_270; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_272 = 10'h110 == io_addr ? 32'h0 : _GEN_271; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_273 = 10'h111 == io_addr ? 32'h0 : _GEN_272; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_274 = 10'h112 == io_addr ? 32'h0 : _GEN_273; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_275 = 10'h113 == io_addr ? 32'h0 : _GEN_274; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_276 = 10'h114 == io_addr ? 32'h0 : _GEN_275; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_277 = 10'h115 == io_addr ? 32'h0 : _GEN_276; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_278 = 10'h116 == io_addr ? 32'h0 : _GEN_277; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_279 = 10'h117 == io_addr ? 32'h0 : _GEN_278; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_280 = 10'h118 == io_addr ? 32'h0 : _GEN_279; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_281 = 10'h119 == io_addr ? 32'h0 : _GEN_280; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_282 = 10'h11a == io_addr ? 32'h0 : _GEN_281; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_283 = 10'h11b == io_addr ? 32'h0 : _GEN_282; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_284 = 10'h11c == io_addr ? 32'h0 : _GEN_283; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_285 = 10'h11d == io_addr ? 32'h0 : _GEN_284; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_286 = 10'h11e == io_addr ? 32'h0 : _GEN_285; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_287 = 10'h11f == io_addr ? 32'h0 : _GEN_286; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_288 = 10'h120 == io_addr ? 32'h0 : _GEN_287; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_289 = 10'h121 == io_addr ? 32'h0 : _GEN_288; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_290 = 10'h122 == io_addr ? 32'h0 : _GEN_289; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_291 = 10'h123 == io_addr ? 32'h0 : _GEN_290; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_292 = 10'h124 == io_addr ? 32'h0 : _GEN_291; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_293 = 10'h125 == io_addr ? 32'h0 : _GEN_292; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_294 = 10'h126 == io_addr ? 32'h0 : _GEN_293; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_295 = 10'h127 == io_addr ? 32'h0 : _GEN_294; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_296 = 10'h128 == io_addr ? 32'h0 : _GEN_295; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_297 = 10'h129 == io_addr ? 32'h0 : _GEN_296; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_298 = 10'h12a == io_addr ? 32'h0 : _GEN_297; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_299 = 10'h12b == io_addr ? 32'h0 : _GEN_298; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_300 = 10'h12c == io_addr ? 32'h0 : _GEN_299; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_301 = 10'h12d == io_addr ? 32'h0 : _GEN_300; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_302 = 10'h12e == io_addr ? 32'h0 : _GEN_301; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_303 = 10'h12f == io_addr ? 32'h0 : _GEN_302; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_304 = 10'h130 == io_addr ? 32'h0 : _GEN_303; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_305 = 10'h131 == io_addr ? 32'h0 : _GEN_304; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_306 = 10'h132 == io_addr ? 32'h0 : _GEN_305; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_307 = 10'h133 == io_addr ? 32'h0 : _GEN_306; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_308 = 10'h134 == io_addr ? 32'h0 : _GEN_307; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_309 = 10'h135 == io_addr ? 32'h0 : _GEN_308; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_310 = 10'h136 == io_addr ? 32'h0 : _GEN_309; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_311 = 10'h137 == io_addr ? 32'h0 : _GEN_310; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_312 = 10'h138 == io_addr ? 32'h0 : _GEN_311; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_313 = 10'h139 == io_addr ? 32'h0 : _GEN_312; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_314 = 10'h13a == io_addr ? 32'h0 : _GEN_313; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_315 = 10'h13b == io_addr ? 32'h0 : _GEN_314; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_316 = 10'h13c == io_addr ? 32'h0 : _GEN_315; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_317 = 10'h13d == io_addr ? 32'h0 : _GEN_316; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_318 = 10'h13e == io_addr ? 32'h0 : _GEN_317; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_319 = 10'h13f == io_addr ? 32'h0 : _GEN_318; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_320 = 10'h140 == io_addr ? 32'h0 : _GEN_319; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_321 = 10'h141 == io_addr ? 32'h0 : _GEN_320; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_322 = 10'h142 == io_addr ? 32'h0 : _GEN_321; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_323 = 10'h143 == io_addr ? 32'h0 : _GEN_322; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_324 = 10'h144 == io_addr ? 32'h0 : _GEN_323; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_325 = 10'h145 == io_addr ? 32'h0 : _GEN_324; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_326 = 10'h146 == io_addr ? 32'h0 : _GEN_325; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_327 = 10'h147 == io_addr ? 32'h0 : _GEN_326; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_328 = 10'h148 == io_addr ? 32'h0 : _GEN_327; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_329 = 10'h149 == io_addr ? 32'h0 : _GEN_328; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_330 = 10'h14a == io_addr ? 32'h0 : _GEN_329; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_331 = 10'h14b == io_addr ? 32'h0 : _GEN_330; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_332 = 10'h14c == io_addr ? 32'h0 : _GEN_331; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_333 = 10'h14d == io_addr ? 32'h0 : _GEN_332; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_334 = 10'h14e == io_addr ? 32'h0 : _GEN_333; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_335 = 10'h14f == io_addr ? 32'h0 : _GEN_334; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_336 = 10'h150 == io_addr ? 32'h0 : _GEN_335; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_337 = 10'h151 == io_addr ? 32'h0 : _GEN_336; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_338 = 10'h152 == io_addr ? 32'h0 : _GEN_337; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_339 = 10'h153 == io_addr ? 32'h0 : _GEN_338; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_340 = 10'h154 == io_addr ? 32'h0 : _GEN_339; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_341 = 10'h155 == io_addr ? 32'h0 : _GEN_340; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_342 = 10'h156 == io_addr ? 32'h0 : _GEN_341; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_343 = 10'h157 == io_addr ? 32'h0 : _GEN_342; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_344 = 10'h158 == io_addr ? 32'h0 : _GEN_343; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_345 = 10'h159 == io_addr ? 32'h0 : _GEN_344; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_346 = 10'h15a == io_addr ? 32'h0 : _GEN_345; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_347 = 10'h15b == io_addr ? 32'h0 : _GEN_346; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_348 = 10'h15c == io_addr ? 32'h0 : _GEN_347; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_349 = 10'h15d == io_addr ? 32'h0 : _GEN_348; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_350 = 10'h15e == io_addr ? 32'h0 : _GEN_349; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_351 = 10'h15f == io_addr ? 32'h0 : _GEN_350; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_352 = 10'h160 == io_addr ? 32'h0 : _GEN_351; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_353 = 10'h161 == io_addr ? 32'h0 : _GEN_352; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_354 = 10'h162 == io_addr ? 32'h0 : _GEN_353; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_355 = 10'h163 == io_addr ? 32'h0 : _GEN_354; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_356 = 10'h164 == io_addr ? 32'h0 : _GEN_355; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_357 = 10'h165 == io_addr ? 32'h0 : _GEN_356; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_358 = 10'h166 == io_addr ? 32'h0 : _GEN_357; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_359 = 10'h167 == io_addr ? 32'h0 : _GEN_358; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_360 = 10'h168 == io_addr ? 32'h0 : _GEN_359; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_361 = 10'h169 == io_addr ? 32'h0 : _GEN_360; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_362 = 10'h16a == io_addr ? 32'h0 : _GEN_361; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_363 = 10'h16b == io_addr ? 32'h0 : _GEN_362; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_364 = 10'h16c == io_addr ? 32'h0 : _GEN_363; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_365 = 10'h16d == io_addr ? 32'h0 : _GEN_364; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_366 = 10'h16e == io_addr ? 32'h0 : _GEN_365; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_367 = 10'h16f == io_addr ? 32'h0 : _GEN_366; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_368 = 10'h170 == io_addr ? 32'h0 : _GEN_367; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_369 = 10'h171 == io_addr ? 32'h0 : _GEN_368; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_370 = 10'h172 == io_addr ? 32'h0 : _GEN_369; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_371 = 10'h173 == io_addr ? 32'h0 : _GEN_370; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_372 = 10'h174 == io_addr ? 32'h0 : _GEN_371; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_373 = 10'h175 == io_addr ? 32'h0 : _GEN_372; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_374 = 10'h176 == io_addr ? 32'h0 : _GEN_373; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_375 = 10'h177 == io_addr ? 32'h0 : _GEN_374; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_376 = 10'h178 == io_addr ? 32'h0 : _GEN_375; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_377 = 10'h179 == io_addr ? 32'h0 : _GEN_376; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_378 = 10'h17a == io_addr ? 32'h0 : _GEN_377; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_379 = 10'h17b == io_addr ? 32'h0 : _GEN_378; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_380 = 10'h17c == io_addr ? 32'h0 : _GEN_379; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_381 = 10'h17d == io_addr ? 32'h0 : _GEN_380; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_382 = 10'h17e == io_addr ? 32'h0 : _GEN_381; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_383 = 10'h17f == io_addr ? 32'h0 : _GEN_382; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_384 = 10'h180 == io_addr ? 32'h0 : _GEN_383; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_385 = 10'h181 == io_addr ? 32'h0 : _GEN_384; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_386 = 10'h182 == io_addr ? 32'h0 : _GEN_385; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_387 = 10'h183 == io_addr ? 32'h0 : _GEN_386; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_388 = 10'h184 == io_addr ? 32'h0 : _GEN_387; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_389 = 10'h185 == io_addr ? 32'h0 : _GEN_388; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_390 = 10'h186 == io_addr ? 32'h0 : _GEN_389; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_391 = 10'h187 == io_addr ? 32'h0 : _GEN_390; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_392 = 10'h188 == io_addr ? 32'h0 : _GEN_391; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_393 = 10'h189 == io_addr ? 32'h0 : _GEN_392; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_394 = 10'h18a == io_addr ? 32'h0 : _GEN_393; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_395 = 10'h18b == io_addr ? 32'h0 : _GEN_394; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_396 = 10'h18c == io_addr ? 32'h0 : _GEN_395; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_397 = 10'h18d == io_addr ? 32'h0 : _GEN_396; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_398 = 10'h18e == io_addr ? 32'h0 : _GEN_397; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_399 = 10'h18f == io_addr ? 32'h0 : _GEN_398; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_400 = 10'h190 == io_addr ? 32'h0 : _GEN_399; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_401 = 10'h191 == io_addr ? 32'h0 : _GEN_400; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_402 = 10'h192 == io_addr ? 32'h0 : _GEN_401; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_403 = 10'h193 == io_addr ? 32'h0 : _GEN_402; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_404 = 10'h194 == io_addr ? 32'h0 : _GEN_403; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_405 = 10'h195 == io_addr ? 32'h0 : _GEN_404; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_406 = 10'h196 == io_addr ? 32'h0 : _GEN_405; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_407 = 10'h197 == io_addr ? 32'h0 : _GEN_406; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_408 = 10'h198 == io_addr ? 32'h0 : _GEN_407; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_409 = 10'h199 == io_addr ? 32'h0 : _GEN_408; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_410 = 10'h19a == io_addr ? 32'h0 : _GEN_409; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_411 = 10'h19b == io_addr ? 32'h0 : _GEN_410; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_412 = 10'h19c == io_addr ? 32'h0 : _GEN_411; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_413 = 10'h19d == io_addr ? 32'h0 : _GEN_412; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_414 = 10'h19e == io_addr ? 32'h0 : _GEN_413; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_415 = 10'h19f == io_addr ? 32'h0 : _GEN_414; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_416 = 10'h1a0 == io_addr ? 32'h0 : _GEN_415; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_417 = 10'h1a1 == io_addr ? 32'h0 : _GEN_416; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_418 = 10'h1a2 == io_addr ? 32'h0 : _GEN_417; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_419 = 10'h1a3 == io_addr ? 32'h0 : _GEN_418; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_420 = 10'h1a4 == io_addr ? 32'h0 : _GEN_419; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_421 = 10'h1a5 == io_addr ? 32'h0 : _GEN_420; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_422 = 10'h1a6 == io_addr ? 32'h0 : _GEN_421; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_423 = 10'h1a7 == io_addr ? 32'h0 : _GEN_422; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_424 = 10'h1a8 == io_addr ? 32'h0 : _GEN_423; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_425 = 10'h1a9 == io_addr ? 32'h0 : _GEN_424; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_426 = 10'h1aa == io_addr ? 32'h0 : _GEN_425; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_427 = 10'h1ab == io_addr ? 32'h0 : _GEN_426; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_428 = 10'h1ac == io_addr ? 32'h0 : _GEN_427; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_429 = 10'h1ad == io_addr ? 32'h0 : _GEN_428; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_430 = 10'h1ae == io_addr ? 32'h0 : _GEN_429; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_431 = 10'h1af == io_addr ? 32'h0 : _GEN_430; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_432 = 10'h1b0 == io_addr ? 32'h0 : _GEN_431; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_433 = 10'h1b1 == io_addr ? 32'h0 : _GEN_432; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_434 = 10'h1b2 == io_addr ? 32'h0 : _GEN_433; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_435 = 10'h1b3 == io_addr ? 32'h0 : _GEN_434; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_436 = 10'h1b4 == io_addr ? 32'h0 : _GEN_435; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_437 = 10'h1b5 == io_addr ? 32'h0 : _GEN_436; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_438 = 10'h1b6 == io_addr ? 32'h0 : _GEN_437; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_439 = 10'h1b7 == io_addr ? 32'h0 : _GEN_438; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_440 = 10'h1b8 == io_addr ? 32'h0 : _GEN_439; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_441 = 10'h1b9 == io_addr ? 32'h0 : _GEN_440; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_442 = 10'h1ba == io_addr ? 32'h0 : _GEN_441; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_443 = 10'h1bb == io_addr ? 32'h0 : _GEN_442; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_444 = 10'h1bc == io_addr ? 32'h0 : _GEN_443; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_445 = 10'h1bd == io_addr ? 32'h0 : _GEN_444; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_446 = 10'h1be == io_addr ? 32'h0 : _GEN_445; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_447 = 10'h1bf == io_addr ? 32'h0 : _GEN_446; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_448 = 10'h1c0 == io_addr ? 32'h0 : _GEN_447; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_449 = 10'h1c1 == io_addr ? 32'h0 : _GEN_448; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_450 = 10'h1c2 == io_addr ? 32'h0 : _GEN_449; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_451 = 10'h1c3 == io_addr ? 32'h0 : _GEN_450; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_452 = 10'h1c4 == io_addr ? 32'h0 : _GEN_451; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_453 = 10'h1c5 == io_addr ? 32'h0 : _GEN_452; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_454 = 10'h1c6 == io_addr ? 32'h0 : _GEN_453; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_455 = 10'h1c7 == io_addr ? 32'h0 : _GEN_454; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_456 = 10'h1c8 == io_addr ? 32'h0 : _GEN_455; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_457 = 10'h1c9 == io_addr ? 32'h0 : _GEN_456; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_458 = 10'h1ca == io_addr ? 32'h0 : _GEN_457; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_459 = 10'h1cb == io_addr ? 32'h0 : _GEN_458; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_460 = 10'h1cc == io_addr ? 32'h0 : _GEN_459; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_461 = 10'h1cd == io_addr ? 32'h0 : _GEN_460; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_462 = 10'h1ce == io_addr ? 32'h0 : _GEN_461; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_463 = 10'h1cf == io_addr ? 32'h0 : _GEN_462; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_464 = 10'h1d0 == io_addr ? 32'h0 : _GEN_463; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_465 = 10'h1d1 == io_addr ? 32'h0 : _GEN_464; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_466 = 10'h1d2 == io_addr ? 32'h0 : _GEN_465; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_467 = 10'h1d3 == io_addr ? 32'h0 : _GEN_466; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_468 = 10'h1d4 == io_addr ? 32'h0 : _GEN_467; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_469 = 10'h1d5 == io_addr ? 32'h0 : _GEN_468; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_470 = 10'h1d6 == io_addr ? 32'h0 : _GEN_469; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_471 = 10'h1d7 == io_addr ? 32'h0 : _GEN_470; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_472 = 10'h1d8 == io_addr ? 32'h0 : _GEN_471; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_473 = 10'h1d9 == io_addr ? 32'h0 : _GEN_472; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_474 = 10'h1da == io_addr ? 32'h0 : _GEN_473; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_475 = 10'h1db == io_addr ? 32'h0 : _GEN_474; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_476 = 10'h1dc == io_addr ? 32'h0 : _GEN_475; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_477 = 10'h1dd == io_addr ? 32'h0 : _GEN_476; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_478 = 10'h1de == io_addr ? 32'h0 : _GEN_477; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_479 = 10'h1df == io_addr ? 32'h0 : _GEN_478; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_480 = 10'h1e0 == io_addr ? 32'h0 : _GEN_479; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_481 = 10'h1e1 == io_addr ? 32'h0 : _GEN_480; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_482 = 10'h1e2 == io_addr ? 32'h0 : _GEN_481; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_483 = 10'h1e3 == io_addr ? 32'h0 : _GEN_482; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_484 = 10'h1e4 == io_addr ? 32'h0 : _GEN_483; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_485 = 10'h1e5 == io_addr ? 32'h0 : _GEN_484; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_486 = 10'h1e6 == io_addr ? 32'h0 : _GEN_485; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_487 = 10'h1e7 == io_addr ? 32'h0 : _GEN_486; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_488 = 10'h1e8 == io_addr ? 32'h0 : _GEN_487; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_489 = 10'h1e9 == io_addr ? 32'h0 : _GEN_488; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_490 = 10'h1ea == io_addr ? 32'h0 : _GEN_489; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_491 = 10'h1eb == io_addr ? 32'h0 : _GEN_490; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_492 = 10'h1ec == io_addr ? 32'h0 : _GEN_491; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_493 = 10'h1ed == io_addr ? 32'h0 : _GEN_492; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_494 = 10'h1ee == io_addr ? 32'h0 : _GEN_493; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_495 = 10'h1ef == io_addr ? 32'h0 : _GEN_494; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_496 = 10'h1f0 == io_addr ? 32'h0 : _GEN_495; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_497 = 10'h1f1 == io_addr ? 32'h0 : _GEN_496; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_498 = 10'h1f2 == io_addr ? 32'h0 : _GEN_497; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_499 = 10'h1f3 == io_addr ? 32'h0 : _GEN_498; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_500 = 10'h1f4 == io_addr ? 32'h0 : _GEN_499; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_501 = 10'h1f5 == io_addr ? 32'h0 : _GEN_500; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_502 = 10'h1f6 == io_addr ? 32'h0 : _GEN_501; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_503 = 10'h1f7 == io_addr ? 32'h0 : _GEN_502; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_504 = 10'h1f8 == io_addr ? 32'h0 : _GEN_503; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_505 = 10'h1f9 == io_addr ? 32'h0 : _GEN_504; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_506 = 10'h1fa == io_addr ? 32'h0 : _GEN_505; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_507 = 10'h1fb == io_addr ? 32'h0 : _GEN_506; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_508 = 10'h1fc == io_addr ? 32'h0 : _GEN_507; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_509 = 10'h1fd == io_addr ? 32'h0 : _GEN_508; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_510 = 10'h1fe == io_addr ? 32'h0 : _GEN_509; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_511 = 10'h1ff == io_addr ? 32'h0 : _GEN_510; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_512 = 10'h200 == io_addr ? 32'h0 : _GEN_511; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_513 = 10'h201 == io_addr ? 32'h0 : _GEN_512; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_514 = 10'h202 == io_addr ? 32'h0 : _GEN_513; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_515 = 10'h203 == io_addr ? 32'h0 : _GEN_514; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_516 = 10'h204 == io_addr ? 32'h0 : _GEN_515; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_517 = 10'h205 == io_addr ? 32'h0 : _GEN_516; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_518 = 10'h206 == io_addr ? 32'h0 : _GEN_517; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_519 = 10'h207 == io_addr ? 32'h0 : _GEN_518; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_520 = 10'h208 == io_addr ? 32'h0 : _GEN_519; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_521 = 10'h209 == io_addr ? 32'h0 : _GEN_520; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_522 = 10'h20a == io_addr ? 32'h0 : _GEN_521; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_523 = 10'h20b == io_addr ? 32'h0 : _GEN_522; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_524 = 10'h20c == io_addr ? 32'h0 : _GEN_523; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_525 = 10'h20d == io_addr ? 32'h0 : _GEN_524; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_526 = 10'h20e == io_addr ? 32'h0 : _GEN_525; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_527 = 10'h20f == io_addr ? 32'h0 : _GEN_526; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_528 = 10'h210 == io_addr ? 32'h0 : _GEN_527; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_529 = 10'h211 == io_addr ? 32'h0 : _GEN_528; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_530 = 10'h212 == io_addr ? 32'h0 : _GEN_529; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_531 = 10'h213 == io_addr ? 32'h0 : _GEN_530; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_532 = 10'h214 == io_addr ? 32'h0 : _GEN_531; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_533 = 10'h215 == io_addr ? 32'h0 : _GEN_532; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_534 = 10'h216 == io_addr ? 32'h0 : _GEN_533; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_535 = 10'h217 == io_addr ? 32'h0 : _GEN_534; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_536 = 10'h218 == io_addr ? 32'h0 : _GEN_535; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_537 = 10'h219 == io_addr ? 32'h0 : _GEN_536; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_538 = 10'h21a == io_addr ? 32'h0 : _GEN_537; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_539 = 10'h21b == io_addr ? 32'h0 : _GEN_538; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_540 = 10'h21c == io_addr ? 32'h0 : _GEN_539; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_541 = 10'h21d == io_addr ? 32'h0 : _GEN_540; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_542 = 10'h21e == io_addr ? 32'h0 : _GEN_541; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_543 = 10'h21f == io_addr ? 32'h0 : _GEN_542; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_544 = 10'h220 == io_addr ? 32'h0 : _GEN_543; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_545 = 10'h221 == io_addr ? 32'h0 : _GEN_544; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_546 = 10'h222 == io_addr ? 32'h0 : _GEN_545; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_547 = 10'h223 == io_addr ? 32'h0 : _GEN_546; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_548 = 10'h224 == io_addr ? 32'h0 : _GEN_547; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_549 = 10'h225 == io_addr ? 32'h0 : _GEN_548; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_550 = 10'h226 == io_addr ? 32'h0 : _GEN_549; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_551 = 10'h227 == io_addr ? 32'h0 : _GEN_550; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_552 = 10'h228 == io_addr ? 32'h0 : _GEN_551; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_553 = 10'h229 == io_addr ? 32'h0 : _GEN_552; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_554 = 10'h22a == io_addr ? 32'h0 : _GEN_553; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_555 = 10'h22b == io_addr ? 32'h0 : _GEN_554; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_556 = 10'h22c == io_addr ? 32'h0 : _GEN_555; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_557 = 10'h22d == io_addr ? 32'h0 : _GEN_556; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_558 = 10'h22e == io_addr ? 32'h0 : _GEN_557; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_559 = 10'h22f == io_addr ? 32'h0 : _GEN_558; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_560 = 10'h230 == io_addr ? 32'h0 : _GEN_559; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_561 = 10'h231 == io_addr ? 32'h0 : _GEN_560; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_562 = 10'h232 == io_addr ? 32'h0 : _GEN_561; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_563 = 10'h233 == io_addr ? 32'h0 : _GEN_562; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_564 = 10'h234 == io_addr ? 32'h0 : _GEN_563; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_565 = 10'h235 == io_addr ? 32'h0 : _GEN_564; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_566 = 10'h236 == io_addr ? 32'h0 : _GEN_565; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_567 = 10'h237 == io_addr ? 32'h0 : _GEN_566; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_568 = 10'h238 == io_addr ? 32'h0 : _GEN_567; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_569 = 10'h239 == io_addr ? 32'h0 : _GEN_568; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_570 = 10'h23a == io_addr ? 32'h0 : _GEN_569; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_571 = 10'h23b == io_addr ? 32'h0 : _GEN_570; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_572 = 10'h23c == io_addr ? 32'h0 : _GEN_571; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_573 = 10'h23d == io_addr ? 32'h0 : _GEN_572; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_574 = 10'h23e == io_addr ? 32'h0 : _GEN_573; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_575 = 10'h23f == io_addr ? 32'h0 : _GEN_574; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_576 = 10'h240 == io_addr ? 32'h0 : _GEN_575; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_577 = 10'h241 == io_addr ? 32'h0 : _GEN_576; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_578 = 10'h242 == io_addr ? 32'h0 : _GEN_577; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_579 = 10'h243 == io_addr ? 32'h0 : _GEN_578; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_580 = 10'h244 == io_addr ? 32'h0 : _GEN_579; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_581 = 10'h245 == io_addr ? 32'h0 : _GEN_580; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_582 = 10'h246 == io_addr ? 32'h0 : _GEN_581; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_583 = 10'h247 == io_addr ? 32'h0 : _GEN_582; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_584 = 10'h248 == io_addr ? 32'h0 : _GEN_583; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_585 = 10'h249 == io_addr ? 32'h0 : _GEN_584; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_586 = 10'h24a == io_addr ? 32'h0 : _GEN_585; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_587 = 10'h24b == io_addr ? 32'h0 : _GEN_586; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_588 = 10'h24c == io_addr ? 32'h0 : _GEN_587; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_589 = 10'h24d == io_addr ? 32'h0 : _GEN_588; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_590 = 10'h24e == io_addr ? 32'h0 : _GEN_589; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_591 = 10'h24f == io_addr ? 32'h0 : _GEN_590; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_592 = 10'h250 == io_addr ? 32'h0 : _GEN_591; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_593 = 10'h251 == io_addr ? 32'h0 : _GEN_592; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_594 = 10'h252 == io_addr ? 32'h0 : _GEN_593; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_595 = 10'h253 == io_addr ? 32'h0 : _GEN_594; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_596 = 10'h254 == io_addr ? 32'h0 : _GEN_595; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_597 = 10'h255 == io_addr ? 32'h0 : _GEN_596; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_598 = 10'h256 == io_addr ? 32'h0 : _GEN_597; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_599 = 10'h257 == io_addr ? 32'h0 : _GEN_598; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_600 = 10'h258 == io_addr ? 32'h0 : _GEN_599; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_601 = 10'h259 == io_addr ? 32'h0 : _GEN_600; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_602 = 10'h25a == io_addr ? 32'h0 : _GEN_601; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_603 = 10'h25b == io_addr ? 32'h0 : _GEN_602; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_604 = 10'h25c == io_addr ? 32'h0 : _GEN_603; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_605 = 10'h25d == io_addr ? 32'h0 : _GEN_604; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_606 = 10'h25e == io_addr ? 32'h0 : _GEN_605; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_607 = 10'h25f == io_addr ? 32'h0 : _GEN_606; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_608 = 10'h260 == io_addr ? 32'h0 : _GEN_607; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_609 = 10'h261 == io_addr ? 32'h0 : _GEN_608; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_610 = 10'h262 == io_addr ? 32'h0 : _GEN_609; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_611 = 10'h263 == io_addr ? 32'h0 : _GEN_610; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_612 = 10'h264 == io_addr ? 32'h0 : _GEN_611; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_613 = 10'h265 == io_addr ? 32'h0 : _GEN_612; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_614 = 10'h266 == io_addr ? 32'h0 : _GEN_613; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_615 = 10'h267 == io_addr ? 32'h0 : _GEN_614; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_616 = 10'h268 == io_addr ? 32'h0 : _GEN_615; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_617 = 10'h269 == io_addr ? 32'h0 : _GEN_616; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_618 = 10'h26a == io_addr ? 32'h0 : _GEN_617; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_619 = 10'h26b == io_addr ? 32'h0 : _GEN_618; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_620 = 10'h26c == io_addr ? 32'h0 : _GEN_619; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_621 = 10'h26d == io_addr ? 32'h0 : _GEN_620; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_622 = 10'h26e == io_addr ? 32'h0 : _GEN_621; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_623 = 10'h26f == io_addr ? 32'h0 : _GEN_622; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_624 = 10'h270 == io_addr ? 32'h0 : _GEN_623; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_625 = 10'h271 == io_addr ? 32'h0 : _GEN_624; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_626 = 10'h272 == io_addr ? 32'h0 : _GEN_625; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_627 = 10'h273 == io_addr ? 32'h0 : _GEN_626; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_628 = 10'h274 == io_addr ? 32'h0 : _GEN_627; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_629 = 10'h275 == io_addr ? 32'h0 : _GEN_628; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_630 = 10'h276 == io_addr ? 32'h0 : _GEN_629; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_631 = 10'h277 == io_addr ? 32'h0 : _GEN_630; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_632 = 10'h278 == io_addr ? 32'h0 : _GEN_631; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_633 = 10'h279 == io_addr ? 32'h0 : _GEN_632; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_634 = 10'h27a == io_addr ? 32'h0 : _GEN_633; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_635 = 10'h27b == io_addr ? 32'h0 : _GEN_634; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_636 = 10'h27c == io_addr ? 32'h0 : _GEN_635; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_637 = 10'h27d == io_addr ? 32'h0 : _GEN_636; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_638 = 10'h27e == io_addr ? 32'h0 : _GEN_637; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_639 = 10'h27f == io_addr ? 32'h0 : _GEN_638; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_640 = 10'h280 == io_addr ? 32'h0 : _GEN_639; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_641 = 10'h281 == io_addr ? 32'h0 : _GEN_640; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_642 = 10'h282 == io_addr ? 32'h0 : _GEN_641; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_643 = 10'h283 == io_addr ? 32'h0 : _GEN_642; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_644 = 10'h284 == io_addr ? 32'h0 : _GEN_643; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_645 = 10'h285 == io_addr ? 32'h0 : _GEN_644; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_646 = 10'h286 == io_addr ? 32'h0 : _GEN_645; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_647 = 10'h287 == io_addr ? 32'h0 : _GEN_646; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_648 = 10'h288 == io_addr ? 32'h0 : _GEN_647; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_649 = 10'h289 == io_addr ? 32'h0 : _GEN_648; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_650 = 10'h28a == io_addr ? 32'h0 : _GEN_649; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_651 = 10'h28b == io_addr ? 32'h0 : _GEN_650; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_652 = 10'h28c == io_addr ? 32'h0 : _GEN_651; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_653 = 10'h28d == io_addr ? 32'h0 : _GEN_652; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_654 = 10'h28e == io_addr ? 32'h0 : _GEN_653; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_655 = 10'h28f == io_addr ? 32'h0 : _GEN_654; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_656 = 10'h290 == io_addr ? 32'h0 : _GEN_655; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_657 = 10'h291 == io_addr ? 32'h0 : _GEN_656; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_658 = 10'h292 == io_addr ? 32'h0 : _GEN_657; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_659 = 10'h293 == io_addr ? 32'h0 : _GEN_658; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_660 = 10'h294 == io_addr ? 32'h0 : _GEN_659; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_661 = 10'h295 == io_addr ? 32'h0 : _GEN_660; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_662 = 10'h296 == io_addr ? 32'h0 : _GEN_661; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_663 = 10'h297 == io_addr ? 32'h0 : _GEN_662; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_664 = 10'h298 == io_addr ? 32'h0 : _GEN_663; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_665 = 10'h299 == io_addr ? 32'h0 : _GEN_664; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_666 = 10'h29a == io_addr ? 32'h0 : _GEN_665; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_667 = 10'h29b == io_addr ? 32'h0 : _GEN_666; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_668 = 10'h29c == io_addr ? 32'h0 : _GEN_667; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_669 = 10'h29d == io_addr ? 32'h0 : _GEN_668; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_670 = 10'h29e == io_addr ? 32'h0 : _GEN_669; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_671 = 10'h29f == io_addr ? 32'h0 : _GEN_670; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_672 = 10'h2a0 == io_addr ? 32'h0 : _GEN_671; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_673 = 10'h2a1 == io_addr ? 32'h0 : _GEN_672; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_674 = 10'h2a2 == io_addr ? 32'h0 : _GEN_673; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_675 = 10'h2a3 == io_addr ? 32'h0 : _GEN_674; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_676 = 10'h2a4 == io_addr ? 32'h0 : _GEN_675; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_677 = 10'h2a5 == io_addr ? 32'h0 : _GEN_676; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_678 = 10'h2a6 == io_addr ? 32'h0 : _GEN_677; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_679 = 10'h2a7 == io_addr ? 32'h0 : _GEN_678; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_680 = 10'h2a8 == io_addr ? 32'h0 : _GEN_679; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_681 = 10'h2a9 == io_addr ? 32'h0 : _GEN_680; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_682 = 10'h2aa == io_addr ? 32'h0 : _GEN_681; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_683 = 10'h2ab == io_addr ? 32'h0 : _GEN_682; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_684 = 10'h2ac == io_addr ? 32'h0 : _GEN_683; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_685 = 10'h2ad == io_addr ? 32'h0 : _GEN_684; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_686 = 10'h2ae == io_addr ? 32'h0 : _GEN_685; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_687 = 10'h2af == io_addr ? 32'h0 : _GEN_686; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_688 = 10'h2b0 == io_addr ? 32'h0 : _GEN_687; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_689 = 10'h2b1 == io_addr ? 32'h0 : _GEN_688; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_690 = 10'h2b2 == io_addr ? 32'h0 : _GEN_689; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_691 = 10'h2b3 == io_addr ? 32'h0 : _GEN_690; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_692 = 10'h2b4 == io_addr ? 32'h0 : _GEN_691; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_693 = 10'h2b5 == io_addr ? 32'h0 : _GEN_692; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_694 = 10'h2b6 == io_addr ? 32'h0 : _GEN_693; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_695 = 10'h2b7 == io_addr ? 32'h0 : _GEN_694; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_696 = 10'h2b8 == io_addr ? 32'h0 : _GEN_695; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_697 = 10'h2b9 == io_addr ? 32'h0 : _GEN_696; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_698 = 10'h2ba == io_addr ? 32'h0 : _GEN_697; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_699 = 10'h2bb == io_addr ? 32'h0 : _GEN_698; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_700 = 10'h2bc == io_addr ? 32'h0 : _GEN_699; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_701 = 10'h2bd == io_addr ? 32'h0 : _GEN_700; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_702 = 10'h2be == io_addr ? 32'h0 : _GEN_701; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_703 = 10'h2bf == io_addr ? 32'h0 : _GEN_702; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_704 = 10'h2c0 == io_addr ? 32'h0 : _GEN_703; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_705 = 10'h2c1 == io_addr ? 32'h0 : _GEN_704; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_706 = 10'h2c2 == io_addr ? 32'h0 : _GEN_705; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_707 = 10'h2c3 == io_addr ? 32'h0 : _GEN_706; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_708 = 10'h2c4 == io_addr ? 32'h0 : _GEN_707; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_709 = 10'h2c5 == io_addr ? 32'h0 : _GEN_708; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_710 = 10'h2c6 == io_addr ? 32'h0 : _GEN_709; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_711 = 10'h2c7 == io_addr ? 32'h0 : _GEN_710; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_712 = 10'h2c8 == io_addr ? 32'h0 : _GEN_711; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_713 = 10'h2c9 == io_addr ? 32'h0 : _GEN_712; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_714 = 10'h2ca == io_addr ? 32'h0 : _GEN_713; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_715 = 10'h2cb == io_addr ? 32'h0 : _GEN_714; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_716 = 10'h2cc == io_addr ? 32'h0 : _GEN_715; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_717 = 10'h2cd == io_addr ? 32'h0 : _GEN_716; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_718 = 10'h2ce == io_addr ? 32'h0 : _GEN_717; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_719 = 10'h2cf == io_addr ? 32'h0 : _GEN_718; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_720 = 10'h2d0 == io_addr ? 32'h0 : _GEN_719; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_721 = 10'h2d1 == io_addr ? 32'h0 : _GEN_720; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_722 = 10'h2d2 == io_addr ? 32'h0 : _GEN_721; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_723 = 10'h2d3 == io_addr ? 32'h0 : _GEN_722; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_724 = 10'h2d4 == io_addr ? 32'h0 : _GEN_723; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_725 = 10'h2d5 == io_addr ? 32'h0 : _GEN_724; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_726 = 10'h2d6 == io_addr ? 32'h0 : _GEN_725; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_727 = 10'h2d7 == io_addr ? 32'h0 : _GEN_726; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_728 = 10'h2d8 == io_addr ? 32'h0 : _GEN_727; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_729 = 10'h2d9 == io_addr ? 32'h0 : _GEN_728; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_730 = 10'h2da == io_addr ? 32'h0 : _GEN_729; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_731 = 10'h2db == io_addr ? 32'h0 : _GEN_730; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_732 = 10'h2dc == io_addr ? 32'h0 : _GEN_731; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_733 = 10'h2dd == io_addr ? 32'h0 : _GEN_732; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_734 = 10'h2de == io_addr ? 32'h0 : _GEN_733; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_735 = 10'h2df == io_addr ? 32'h0 : _GEN_734; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_736 = 10'h2e0 == io_addr ? 32'h0 : _GEN_735; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_737 = 10'h2e1 == io_addr ? 32'h0 : _GEN_736; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_738 = 10'h2e2 == io_addr ? 32'h0 : _GEN_737; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_739 = 10'h2e3 == io_addr ? 32'h0 : _GEN_738; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_740 = 10'h2e4 == io_addr ? 32'h0 : _GEN_739; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_741 = 10'h2e5 == io_addr ? 32'h0 : _GEN_740; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_742 = 10'h2e6 == io_addr ? 32'h0 : _GEN_741; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_743 = 10'h2e7 == io_addr ? 32'h0 : _GEN_742; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_744 = 10'h2e8 == io_addr ? 32'h0 : _GEN_743; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_745 = 10'h2e9 == io_addr ? 32'h0 : _GEN_744; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_746 = 10'h2ea == io_addr ? 32'h0 : _GEN_745; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_747 = 10'h2eb == io_addr ? 32'h0 : _GEN_746; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_748 = 10'h2ec == io_addr ? 32'h0 : _GEN_747; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_749 = 10'h2ed == io_addr ? 32'h0 : _GEN_748; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_750 = 10'h2ee == io_addr ? 32'h0 : _GEN_749; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_751 = 10'h2ef == io_addr ? 32'h0 : _GEN_750; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_752 = 10'h2f0 == io_addr ? 32'h0 : _GEN_751; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_753 = 10'h2f1 == io_addr ? 32'h0 : _GEN_752; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_754 = 10'h2f2 == io_addr ? 32'h0 : _GEN_753; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_755 = 10'h2f3 == io_addr ? 32'h0 : _GEN_754; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_756 = 10'h2f4 == io_addr ? 32'h0 : _GEN_755; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_757 = 10'h2f5 == io_addr ? 32'h0 : _GEN_756; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_758 = 10'h2f6 == io_addr ? 32'h0 : _GEN_757; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_759 = 10'h2f7 == io_addr ? 32'h0 : _GEN_758; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_760 = 10'h2f8 == io_addr ? 32'h0 : _GEN_759; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_761 = 10'h2f9 == io_addr ? 32'h0 : _GEN_760; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_762 = 10'h2fa == io_addr ? 32'h0 : _GEN_761; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_763 = 10'h2fb == io_addr ? 32'h0 : _GEN_762; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_764 = 10'h2fc == io_addr ? 32'h0 : _GEN_763; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_765 = 10'h2fd == io_addr ? 32'h0 : _GEN_764; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_766 = 10'h2fe == io_addr ? 32'h0 : _GEN_765; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_767 = 10'h2ff == io_addr ? 32'h0 : _GEN_766; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_768 = 10'h300 == io_addr ? 32'h0 : _GEN_767; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_769 = 10'h301 == io_addr ? 32'h0 : _GEN_768; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_770 = 10'h302 == io_addr ? 32'h0 : _GEN_769; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_771 = 10'h303 == io_addr ? 32'h0 : _GEN_770; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_772 = 10'h304 == io_addr ? 32'h0 : _GEN_771; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_773 = 10'h305 == io_addr ? 32'h0 : _GEN_772; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_774 = 10'h306 == io_addr ? 32'h0 : _GEN_773; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_775 = 10'h307 == io_addr ? 32'h0 : _GEN_774; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_776 = 10'h308 == io_addr ? 32'h0 : _GEN_775; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_777 = 10'h309 == io_addr ? 32'h0 : _GEN_776; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_778 = 10'h30a == io_addr ? 32'h0 : _GEN_777; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_779 = 10'h30b == io_addr ? 32'h0 : _GEN_778; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_780 = 10'h30c == io_addr ? 32'h0 : _GEN_779; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_781 = 10'h30d == io_addr ? 32'h0 : _GEN_780; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_782 = 10'h30e == io_addr ? 32'h0 : _GEN_781; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_783 = 10'h30f == io_addr ? 32'h0 : _GEN_782; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_784 = 10'h310 == io_addr ? 32'h0 : _GEN_783; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_785 = 10'h311 == io_addr ? 32'h0 : _GEN_784; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_786 = 10'h312 == io_addr ? 32'h0 : _GEN_785; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_787 = 10'h313 == io_addr ? 32'h0 : _GEN_786; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_788 = 10'h314 == io_addr ? 32'h0 : _GEN_787; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_789 = 10'h315 == io_addr ? 32'h0 : _GEN_788; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_790 = 10'h316 == io_addr ? 32'h0 : _GEN_789; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_791 = 10'h317 == io_addr ? 32'h0 : _GEN_790; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_792 = 10'h318 == io_addr ? 32'h0 : _GEN_791; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_793 = 10'h319 == io_addr ? 32'h0 : _GEN_792; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_794 = 10'h31a == io_addr ? 32'h0 : _GEN_793; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_795 = 10'h31b == io_addr ? 32'h0 : _GEN_794; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_796 = 10'h31c == io_addr ? 32'h0 : _GEN_795; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_797 = 10'h31d == io_addr ? 32'h0 : _GEN_796; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_798 = 10'h31e == io_addr ? 32'h0 : _GEN_797; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_799 = 10'h31f == io_addr ? 32'h0 : _GEN_798; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_800 = 10'h320 == io_addr ? 32'h0 : _GEN_799; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_801 = 10'h321 == io_addr ? 32'h0 : _GEN_800; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_802 = 10'h322 == io_addr ? 32'h0 : _GEN_801; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_803 = 10'h323 == io_addr ? 32'h0 : _GEN_802; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_804 = 10'h324 == io_addr ? 32'h0 : _GEN_803; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_805 = 10'h325 == io_addr ? 32'h0 : _GEN_804; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_806 = 10'h326 == io_addr ? 32'h0 : _GEN_805; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_807 = 10'h327 == io_addr ? 32'h0 : _GEN_806; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_808 = 10'h328 == io_addr ? 32'h0 : _GEN_807; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_809 = 10'h329 == io_addr ? 32'h0 : _GEN_808; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_810 = 10'h32a == io_addr ? 32'h0 : _GEN_809; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_811 = 10'h32b == io_addr ? 32'h0 : _GEN_810; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_812 = 10'h32c == io_addr ? 32'h0 : _GEN_811; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_813 = 10'h32d == io_addr ? 32'h0 : _GEN_812; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_814 = 10'h32e == io_addr ? 32'h0 : _GEN_813; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_815 = 10'h32f == io_addr ? 32'h0 : _GEN_814; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_816 = 10'h330 == io_addr ? 32'h0 : _GEN_815; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_817 = 10'h331 == io_addr ? 32'h0 : _GEN_816; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_818 = 10'h332 == io_addr ? 32'h0 : _GEN_817; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_819 = 10'h333 == io_addr ? 32'h0 : _GEN_818; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_820 = 10'h334 == io_addr ? 32'h0 : _GEN_819; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_821 = 10'h335 == io_addr ? 32'h0 : _GEN_820; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_822 = 10'h336 == io_addr ? 32'h0 : _GEN_821; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_823 = 10'h337 == io_addr ? 32'h0 : _GEN_822; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_824 = 10'h338 == io_addr ? 32'h0 : _GEN_823; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_825 = 10'h339 == io_addr ? 32'h0 : _GEN_824; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_826 = 10'h33a == io_addr ? 32'h0 : _GEN_825; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_827 = 10'h33b == io_addr ? 32'h0 : _GEN_826; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_828 = 10'h33c == io_addr ? 32'h0 : _GEN_827; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_829 = 10'h33d == io_addr ? 32'h0 : _GEN_828; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_830 = 10'h33e == io_addr ? 32'h0 : _GEN_829; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_831 = 10'h33f == io_addr ? 32'h0 : _GEN_830; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_832 = 10'h340 == io_addr ? 32'h0 : _GEN_831; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_833 = 10'h341 == io_addr ? 32'h0 : _GEN_832; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_834 = 10'h342 == io_addr ? 32'h0 : _GEN_833; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_835 = 10'h343 == io_addr ? 32'h0 : _GEN_834; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_836 = 10'h344 == io_addr ? 32'h0 : _GEN_835; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_837 = 10'h345 == io_addr ? 32'h0 : _GEN_836; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_838 = 10'h346 == io_addr ? 32'h0 : _GEN_837; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_839 = 10'h347 == io_addr ? 32'h0 : _GEN_838; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_840 = 10'h348 == io_addr ? 32'h0 : _GEN_839; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_841 = 10'h349 == io_addr ? 32'h0 : _GEN_840; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_842 = 10'h34a == io_addr ? 32'h0 : _GEN_841; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_843 = 10'h34b == io_addr ? 32'h0 : _GEN_842; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_844 = 10'h34c == io_addr ? 32'h0 : _GEN_843; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_845 = 10'h34d == io_addr ? 32'h0 : _GEN_844; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_846 = 10'h34e == io_addr ? 32'h0 : _GEN_845; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_847 = 10'h34f == io_addr ? 32'h0 : _GEN_846; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_848 = 10'h350 == io_addr ? 32'h0 : _GEN_847; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_849 = 10'h351 == io_addr ? 32'h0 : _GEN_848; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_850 = 10'h352 == io_addr ? 32'h0 : _GEN_849; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_851 = 10'h353 == io_addr ? 32'h0 : _GEN_850; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_852 = 10'h354 == io_addr ? 32'h0 : _GEN_851; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_853 = 10'h355 == io_addr ? 32'h0 : _GEN_852; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_854 = 10'h356 == io_addr ? 32'h0 : _GEN_853; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_855 = 10'h357 == io_addr ? 32'h0 : _GEN_854; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_856 = 10'h358 == io_addr ? 32'h0 : _GEN_855; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_857 = 10'h359 == io_addr ? 32'h0 : _GEN_856; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_858 = 10'h35a == io_addr ? 32'h0 : _GEN_857; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_859 = 10'h35b == io_addr ? 32'h0 : _GEN_858; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_860 = 10'h35c == io_addr ? 32'h0 : _GEN_859; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_861 = 10'h35d == io_addr ? 32'h0 : _GEN_860; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_862 = 10'h35e == io_addr ? 32'h0 : _GEN_861; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_863 = 10'h35f == io_addr ? 32'h0 : _GEN_862; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_864 = 10'h360 == io_addr ? 32'h0 : _GEN_863; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_865 = 10'h361 == io_addr ? 32'h0 : _GEN_864; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_866 = 10'h362 == io_addr ? 32'h0 : _GEN_865; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_867 = 10'h363 == io_addr ? 32'h0 : _GEN_866; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_868 = 10'h364 == io_addr ? 32'h0 : _GEN_867; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_869 = 10'h365 == io_addr ? 32'h0 : _GEN_868; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_870 = 10'h366 == io_addr ? 32'h0 : _GEN_869; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_871 = 10'h367 == io_addr ? 32'h0 : _GEN_870; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_872 = 10'h368 == io_addr ? 32'h0 : _GEN_871; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_873 = 10'h369 == io_addr ? 32'h0 : _GEN_872; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_874 = 10'h36a == io_addr ? 32'h0 : _GEN_873; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_875 = 10'h36b == io_addr ? 32'h0 : _GEN_874; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_876 = 10'h36c == io_addr ? 32'h0 : _GEN_875; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_877 = 10'h36d == io_addr ? 32'h0 : _GEN_876; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_878 = 10'h36e == io_addr ? 32'h0 : _GEN_877; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_879 = 10'h36f == io_addr ? 32'h0 : _GEN_878; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_880 = 10'h370 == io_addr ? 32'h0 : _GEN_879; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_881 = 10'h371 == io_addr ? 32'h0 : _GEN_880; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_882 = 10'h372 == io_addr ? 32'h0 : _GEN_881; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_883 = 10'h373 == io_addr ? 32'h0 : _GEN_882; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_884 = 10'h374 == io_addr ? 32'h0 : _GEN_883; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_885 = 10'h375 == io_addr ? 32'h0 : _GEN_884; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_886 = 10'h376 == io_addr ? 32'h0 : _GEN_885; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_887 = 10'h377 == io_addr ? 32'h0 : _GEN_886; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_888 = 10'h378 == io_addr ? 32'h0 : _GEN_887; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_889 = 10'h379 == io_addr ? 32'h0 : _GEN_888; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_890 = 10'h37a == io_addr ? 32'h0 : _GEN_889; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_891 = 10'h37b == io_addr ? 32'h0 : _GEN_890; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_892 = 10'h37c == io_addr ? 32'h0 : _GEN_891; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_893 = 10'h37d == io_addr ? 32'h0 : _GEN_892; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_894 = 10'h37e == io_addr ? 32'h0 : _GEN_893; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_895 = 10'h37f == io_addr ? 32'h0 : _GEN_894; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_896 = 10'h380 == io_addr ? 32'h0 : _GEN_895; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_897 = 10'h381 == io_addr ? 32'h0 : _GEN_896; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_898 = 10'h382 == io_addr ? 32'h0 : _GEN_897; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_899 = 10'h383 == io_addr ? 32'h0 : _GEN_898; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_900 = 10'h384 == io_addr ? 32'h0 : _GEN_899; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_901 = 10'h385 == io_addr ? 32'h0 : _GEN_900; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_902 = 10'h386 == io_addr ? 32'h0 : _GEN_901; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_903 = 10'h387 == io_addr ? 32'h0 : _GEN_902; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_904 = 10'h388 == io_addr ? 32'h0 : _GEN_903; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_905 = 10'h389 == io_addr ? 32'h0 : _GEN_904; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_906 = 10'h38a == io_addr ? 32'h0 : _GEN_905; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_907 = 10'h38b == io_addr ? 32'h0 : _GEN_906; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_908 = 10'h38c == io_addr ? 32'h0 : _GEN_907; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_909 = 10'h38d == io_addr ? 32'h0 : _GEN_908; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_910 = 10'h38e == io_addr ? 32'h0 : _GEN_909; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_911 = 10'h38f == io_addr ? 32'h0 : _GEN_910; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_912 = 10'h390 == io_addr ? 32'h0 : _GEN_911; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_913 = 10'h391 == io_addr ? 32'h0 : _GEN_912; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_914 = 10'h392 == io_addr ? 32'h0 : _GEN_913; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_915 = 10'h393 == io_addr ? 32'h0 : _GEN_914; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_916 = 10'h394 == io_addr ? 32'h0 : _GEN_915; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_917 = 10'h395 == io_addr ? 32'h0 : _GEN_916; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_918 = 10'h396 == io_addr ? 32'h0 : _GEN_917; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_919 = 10'h397 == io_addr ? 32'h0 : _GEN_918; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_920 = 10'h398 == io_addr ? 32'h0 : _GEN_919; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_921 = 10'h399 == io_addr ? 32'h0 : _GEN_920; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_922 = 10'h39a == io_addr ? 32'h0 : _GEN_921; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_923 = 10'h39b == io_addr ? 32'h0 : _GEN_922; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_924 = 10'h39c == io_addr ? 32'h0 : _GEN_923; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_925 = 10'h39d == io_addr ? 32'h0 : _GEN_924; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_926 = 10'h39e == io_addr ? 32'h0 : _GEN_925; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_927 = 10'h39f == io_addr ? 32'h0 : _GEN_926; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_928 = 10'h3a0 == io_addr ? 32'h0 : _GEN_927; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_929 = 10'h3a1 == io_addr ? 32'h0 : _GEN_928; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_930 = 10'h3a2 == io_addr ? 32'h0 : _GEN_929; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_931 = 10'h3a3 == io_addr ? 32'h0 : _GEN_930; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_932 = 10'h3a4 == io_addr ? 32'h0 : _GEN_931; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_933 = 10'h3a5 == io_addr ? 32'h0 : _GEN_932; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_934 = 10'h3a6 == io_addr ? 32'h0 : _GEN_933; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_935 = 10'h3a7 == io_addr ? 32'h0 : _GEN_934; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_936 = 10'h3a8 == io_addr ? 32'h0 : _GEN_935; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_937 = 10'h3a9 == io_addr ? 32'h0 : _GEN_936; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_938 = 10'h3aa == io_addr ? 32'h0 : _GEN_937; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_939 = 10'h3ab == io_addr ? 32'h0 : _GEN_938; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_940 = 10'h3ac == io_addr ? 32'h0 : _GEN_939; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_941 = 10'h3ad == io_addr ? 32'h0 : _GEN_940; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_942 = 10'h3ae == io_addr ? 32'h0 : _GEN_941; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_943 = 10'h3af == io_addr ? 32'h0 : _GEN_942; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_944 = 10'h3b0 == io_addr ? 32'h0 : _GEN_943; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_945 = 10'h3b1 == io_addr ? 32'h0 : _GEN_944; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_946 = 10'h3b2 == io_addr ? 32'h0 : _GEN_945; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_947 = 10'h3b3 == io_addr ? 32'h0 : _GEN_946; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_948 = 10'h3b4 == io_addr ? 32'h0 : _GEN_947; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_949 = 10'h3b5 == io_addr ? 32'h0 : _GEN_948; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_950 = 10'h3b6 == io_addr ? 32'h0 : _GEN_949; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_951 = 10'h3b7 == io_addr ? 32'h0 : _GEN_950; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_952 = 10'h3b8 == io_addr ? 32'h0 : _GEN_951; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_953 = 10'h3b9 == io_addr ? 32'h0 : _GEN_952; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_954 = 10'h3ba == io_addr ? 32'h0 : _GEN_953; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_955 = 10'h3bb == io_addr ? 32'h0 : _GEN_954; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_956 = 10'h3bc == io_addr ? 32'h0 : _GEN_955; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_957 = 10'h3bd == io_addr ? 32'h0 : _GEN_956; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_958 = 10'h3be == io_addr ? 32'h0 : _GEN_957; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_959 = 10'h3bf == io_addr ? 32'h0 : _GEN_958; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_960 = 10'h3c0 == io_addr ? 32'h0 : _GEN_959; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_961 = 10'h3c1 == io_addr ? 32'h0 : _GEN_960; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_962 = 10'h3c2 == io_addr ? 32'h0 : _GEN_961; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_963 = 10'h3c3 == io_addr ? 32'h0 : _GEN_962; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_964 = 10'h3c4 == io_addr ? 32'h0 : _GEN_963; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_965 = 10'h3c5 == io_addr ? 32'h0 : _GEN_964; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_966 = 10'h3c6 == io_addr ? 32'h0 : _GEN_965; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_967 = 10'h3c7 == io_addr ? 32'h0 : _GEN_966; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_968 = 10'h3c8 == io_addr ? 32'h0 : _GEN_967; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_969 = 10'h3c9 == io_addr ? 32'h0 : _GEN_968; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_970 = 10'h3ca == io_addr ? 32'h0 : _GEN_969; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_971 = 10'h3cb == io_addr ? 32'h0 : _GEN_970; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_972 = 10'h3cc == io_addr ? 32'h0 : _GEN_971; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_973 = 10'h3cd == io_addr ? 32'h0 : _GEN_972; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_974 = 10'h3ce == io_addr ? 32'h0 : _GEN_973; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_975 = 10'h3cf == io_addr ? 32'h0 : _GEN_974; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_976 = 10'h3d0 == io_addr ? 32'h0 : _GEN_975; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_977 = 10'h3d1 == io_addr ? 32'h0 : _GEN_976; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_978 = 10'h3d2 == io_addr ? 32'h0 : _GEN_977; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_979 = 10'h3d3 == io_addr ? 32'h0 : _GEN_978; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_980 = 10'h3d4 == io_addr ? 32'h0 : _GEN_979; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_981 = 10'h3d5 == io_addr ? 32'h0 : _GEN_980; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_982 = 10'h3d6 == io_addr ? 32'h0 : _GEN_981; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_983 = 10'h3d7 == io_addr ? 32'h0 : _GEN_982; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_984 = 10'h3d8 == io_addr ? 32'h0 : _GEN_983; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_985 = 10'h3d9 == io_addr ? 32'h0 : _GEN_984; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_986 = 10'h3da == io_addr ? 32'h0 : _GEN_985; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_987 = 10'h3db == io_addr ? 32'h0 : _GEN_986; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_988 = 10'h3dc == io_addr ? 32'h0 : _GEN_987; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_989 = 10'h3dd == io_addr ? 32'h0 : _GEN_988; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_990 = 10'h3de == io_addr ? 32'h0 : _GEN_989; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_991 = 10'h3df == io_addr ? 32'h0 : _GEN_990; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_992 = 10'h3e0 == io_addr ? 32'h0 : _GEN_991; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_993 = 10'h3e1 == io_addr ? 32'h0 : _GEN_992; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_994 = 10'h3e2 == io_addr ? 32'h0 : _GEN_993; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_995 = 10'h3e3 == io_addr ? 32'h0 : _GEN_994; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_996 = 10'h3e4 == io_addr ? 32'h0 : _GEN_995; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_997 = 10'h3e5 == io_addr ? 32'h0 : _GEN_996; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_998 = 10'h3e6 == io_addr ? 32'h0 : _GEN_997; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_999 = 10'h3e7 == io_addr ? 32'h0 : _GEN_998; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1000 = 10'h3e8 == io_addr ? 32'h0 : _GEN_999; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1001 = 10'h3e9 == io_addr ? 32'h0 : _GEN_1000; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1002 = 10'h3ea == io_addr ? 32'h0 : _GEN_1001; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1003 = 10'h3eb == io_addr ? 32'h0 : _GEN_1002; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1004 = 10'h3ec == io_addr ? 32'h0 : _GEN_1003; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1005 = 10'h3ed == io_addr ? 32'h0 : _GEN_1004; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1006 = 10'h3ee == io_addr ? 32'h0 : _GEN_1005; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1007 = 10'h3ef == io_addr ? 32'h0 : _GEN_1006; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1008 = 10'h3f0 == io_addr ? 32'h0 : _GEN_1007; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1009 = 10'h3f1 == io_addr ? 32'h0 : _GEN_1008; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1010 = 10'h3f2 == io_addr ? 32'h0 : _GEN_1009; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1011 = 10'h3f3 == io_addr ? 32'h0 : _GEN_1010; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1012 = 10'h3f4 == io_addr ? 32'h0 : _GEN_1011; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1013 = 10'h3f5 == io_addr ? 32'h0 : _GEN_1012; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1014 = 10'h3f6 == io_addr ? 32'h0 : _GEN_1013; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1015 = 10'h3f7 == io_addr ? 32'h0 : _GEN_1014; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1016 = 10'h3f8 == io_addr ? 32'h0 : _GEN_1015; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1017 = 10'h3f9 == io_addr ? 32'h0 : _GEN_1016; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1018 = 10'h3fa == io_addr ? 32'h0 : _GEN_1017; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1019 = 10'h3fb == io_addr ? 32'h0 : _GEN_1018; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1020 = 10'h3fc == io_addr ? 32'h0 : _GEN_1019; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1021 = 10'h3fd == io_addr ? 32'h0 : _GEN_1020; // @[InstrMemoryTest.scala 20:{24,24}]
  wire [31:0] _GEN_1022 = 10'h3fe == io_addr ? 32'h0 : _GEN_1021; // @[InstrMemoryTest.scala 20:{24,24}]
  assign io_dataOut = 10'h3ff == io_addr ? 32'h0 : _GEN_1022; // @[InstrMemoryTest.scala 20:{24,24}]
  always @(posedge clock) begin
    if (reset) begin // @[InstrMemoryTest.scala 20:24]
      dataReg <= 32'h0; // @[InstrMemoryTest.scala 20:24]
    end else if (10'h3ff == io_addr) begin // @[InstrMemoryTest.scala 20:24]
      dataReg <= 32'h0; // @[InstrMemoryTest.scala 20:24]
    end else if (10'h3fe == io_addr) begin // @[InstrMemoryTest.scala 20:24]
      dataReg <= 32'h0; // @[InstrMemoryTest.scala 20:24]
    end else if (10'h3fd == io_addr) begin // @[InstrMemoryTest.scala 20:24]
      dataReg <= 32'h0; // @[InstrMemoryTest.scala 20:24]
    end else begin
      dataReg <= _GEN_1020;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dataReg = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFStage(
  input         clock,
  input         reset,
  output [31:0] io_instruction
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  instrMem_clock; // @[IFStage.scala 24:24]
  wire  instrMem_reset; // @[IFStage.scala 24:24]
  wire [9:0] instrMem_io_addr; // @[IFStage.scala 24:24]
  wire [31:0] instrMem_io_dataOut; // @[IFStage.scala 24:24]
  reg [31:0] PC; // @[IFStage.scala 18:19]
  wire [31:0] NextInstrAdd = PC + 32'h4; // @[IFStage.scala 19:74]
  wire [31:0] _instrMem_io_addr_T = {{2'd0}, NextInstrAdd[31:2]}; // @[IFStage.scala 26:36]
  InstrMemoryTest instrMem ( // @[IFStage.scala 24:24]
    .clock(instrMem_clock),
    .reset(instrMem_reset),
    .io_addr(instrMem_io_addr),
    .io_dataOut(instrMem_io_dataOut)
  );
  assign io_instruction = instrMem_io_dataOut; // @[IFStage.scala 27:18]
  assign instrMem_clock = clock;
  assign instrMem_reset = reset;
  assign instrMem_io_addr = _instrMem_io_addr_T[9:0]; // @[IFStage.scala 26:20]
  always @(posedge clock) begin
    if (reset) begin // @[IFStage.scala 18:19]
      PC <= 32'hfffffffc; // @[IFStage.scala 18:19]
    end else begin
      PC <= NextInstrAdd; // @[IFStage.scala 21:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  PC = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstructionDecoder(
  input  [31:0] io_instruction,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [2:0]  io_funct3,
  output [6:0]  io_funct7,
  output [2:0]  io_instrType,
  output [6:0]  io_opcode
);
  wire [2:0] _GEN_0 = 7'h37 == io_opcode ? 3'h4 : 3'h0; // @[IDStage.scala 27:16 30:21 56:20]
  wire [2:0] _GEN_1 = 7'h17 == io_opcode ? 3'h4 : _GEN_0; // @[IDStage.scala 30:21 53:20]
  wire [2:0] _GEN_2 = 7'h67 == io_opcode ? 3'h1 : _GEN_1; // @[IDStage.scala 30:21 50:20]
  wire [2:0] _GEN_3 = 7'h6f == io_opcode ? 3'h5 : _GEN_2; // @[IDStage.scala 30:21 47:20]
  wire [2:0] _GEN_4 = 7'h63 == io_opcode ? 3'h3 : _GEN_3; // @[IDStage.scala 30:21 44:20]
  wire [2:0] _GEN_5 = 7'h23 == io_opcode ? 3'h2 : _GEN_4; // @[IDStage.scala 30:21 41:20]
  wire [2:0] _GEN_6 = 7'h3 == io_opcode ? 3'h1 : _GEN_5; // @[IDStage.scala 30:21 38:20]
  wire [2:0] _GEN_7 = 7'h13 == io_opcode ? 3'h1 : _GEN_6; // @[IDStage.scala 30:21 35:20]
  wire [6:0] _GEN_9 = io_funct3 == 3'h1 | io_funct3 == 3'h5 | io_funct3 == 3'h5 ? io_instruction[31:25] : 7'h0; // @[IDStage.scala 72:108 26:13 74:19]
  wire [4:0] _GEN_10 = 3'h4 == io_instrType ? io_instruction[11:7] : 5'h0; // @[IDStage.scala 60:24 91:13 24:9]
  wire [4:0] _GEN_11 = 3'h5 == io_instrType ? io_instruction[11:7] : _GEN_10; // @[IDStage.scala 60:24 88:13]
  wire [4:0] _GEN_12 = 3'h3 == io_instrType ? io_instruction[19:15] : 5'h0; // @[IDStage.scala 22:10 60:24 83:14]
  wire [4:0] _GEN_13 = 3'h3 == io_instrType ? io_instruction[24:20] : 5'h0; // @[IDStage.scala 23:10 60:24 84:14]
  wire [2:0] _GEN_14 = 3'h3 == io_instrType ? io_instruction[14:12] : 3'h0; // @[IDStage.scala 25:13 60:24 85:17]
  wire [4:0] _GEN_15 = 3'h3 == io_instrType ? 5'h0 : _GEN_11; // @[IDStage.scala 60:24 24:9]
  wire [4:0] _GEN_16 = 3'h2 == io_instrType ? io_instruction[19:15] : _GEN_12; // @[IDStage.scala 60:24 78:14]
  wire [4:0] _GEN_17 = 3'h2 == io_instrType ? io_instruction[24:20] : _GEN_13; // @[IDStage.scala 60:24 79:14]
  wire [2:0] _GEN_18 = 3'h2 == io_instrType ? io_instruction[14:12] : _GEN_14; // @[IDStage.scala 60:24 80:17]
  wire [4:0] _GEN_19 = 3'h2 == io_instrType ? 5'h0 : _GEN_15; // @[IDStage.scala 60:24 24:9]
  wire [4:0] _GEN_20 = 3'h1 == io_instrType ? io_instruction[19:15] : _GEN_16; // @[IDStage.scala 60:24 69:14]
  wire [2:0] _GEN_21 = 3'h1 == io_instrType ? io_instruction[14:12] : _GEN_18; // @[IDStage.scala 60:24 70:17]
  wire [4:0] _GEN_22 = 3'h1 == io_instrType ? io_instruction[11:7] : _GEN_19; // @[IDStage.scala 60:24 71:13]
  wire [6:0] _GEN_23 = 3'h1 == io_instrType ? _GEN_9 : 7'h0; // @[IDStage.scala 26:13 60:24]
  wire [4:0] _GEN_24 = 3'h1 == io_instrType ? 5'h0 : _GEN_17; // @[IDStage.scala 23:10 60:24]
  assign io_rs1 = 3'h0 == io_instrType ? io_instruction[19:15] : _GEN_20; // @[IDStage.scala 60:24 62:14]
  assign io_rs2 = 3'h0 == io_instrType ? io_instruction[24:20] : _GEN_24; // @[IDStage.scala 60:24 63:14]
  assign io_rd = 3'h0 == io_instrType ? io_instruction[11:7] : _GEN_22; // @[IDStage.scala 60:24 64:13]
  assign io_funct3 = 3'h0 == io_instrType ? io_instruction[14:12] : _GEN_21; // @[IDStage.scala 60:24 65:17]
  assign io_funct7 = 3'h0 == io_instrType ? io_instruction[31:25] : _GEN_23; // @[IDStage.scala 60:24 66:17]
  assign io_instrType = 7'h33 == io_opcode ? 3'h0 : _GEN_7; // @[IDStage.scala 30:21 32:20]
  assign io_opcode = io_instruction[6:0]; // @[IDStage.scala 28:30]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [31:0] io_writeData,
  input  [4:0]  io_rd,
  input         io_writeEnable,
  output [31:0] io_operand1,
  output [31:0] io_operand2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] RegFile_0; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_1; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_2; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_3; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_4; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_5; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_6; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_7; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_8; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_9; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_10; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_11; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_12; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_13; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_14; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_15; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_16; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_17; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_18; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_19; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_20; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_21; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_22; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_23; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_24; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_25; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_26; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_27; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_28; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_29; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_30; // @[RegisterFile.scala 19:25]
  reg [31:0] RegFile_31; // @[RegisterFile.scala 19:25]
  wire [31:0] _GEN_0 = 5'h0 == io_rd ? io_writeData : RegFile_0; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_1 = 5'h1 == io_rd ? io_writeData : RegFile_1; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_2 = 5'h2 == io_rd ? io_writeData : RegFile_2; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_3 = 5'h3 == io_rd ? io_writeData : RegFile_3; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_4 = 5'h4 == io_rd ? io_writeData : RegFile_4; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_5 = 5'h5 == io_rd ? io_writeData : RegFile_5; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_6 = 5'h6 == io_rd ? io_writeData : RegFile_6; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_7 = 5'h7 == io_rd ? io_writeData : RegFile_7; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_8 = 5'h8 == io_rd ? io_writeData : RegFile_8; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_9 = 5'h9 == io_rd ? io_writeData : RegFile_9; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_10 = 5'ha == io_rd ? io_writeData : RegFile_10; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_11 = 5'hb == io_rd ? io_writeData : RegFile_11; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_12 = 5'hc == io_rd ? io_writeData : RegFile_12; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_13 = 5'hd == io_rd ? io_writeData : RegFile_13; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_14 = 5'he == io_rd ? io_writeData : RegFile_14; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_15 = 5'hf == io_rd ? io_writeData : RegFile_15; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_16 = 5'h10 == io_rd ? io_writeData : RegFile_16; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_17 = 5'h11 == io_rd ? io_writeData : RegFile_17; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_18 = 5'h12 == io_rd ? io_writeData : RegFile_18; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_19 = 5'h13 == io_rd ? io_writeData : RegFile_19; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_20 = 5'h14 == io_rd ? io_writeData : RegFile_20; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_21 = 5'h15 == io_rd ? io_writeData : RegFile_21; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_22 = 5'h16 == io_rd ? io_writeData : RegFile_22; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_23 = 5'h17 == io_rd ? io_writeData : RegFile_23; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_24 = 5'h18 == io_rd ? io_writeData : RegFile_24; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_25 = 5'h19 == io_rd ? io_writeData : RegFile_25; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_26 = 5'h1a == io_rd ? io_writeData : RegFile_26; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_27 = 5'h1b == io_rd ? io_writeData : RegFile_27; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_28 = 5'h1c == io_rd ? io_writeData : RegFile_28; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_29 = 5'h1d == io_rd ? io_writeData : RegFile_29; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_30 = 5'h1e == io_rd ? io_writeData : RegFile_30; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire [31:0] _GEN_31 = 5'h1f == io_rd ? io_writeData : RegFile_31; // @[RegisterFile.scala 26:{20,20} 19:25]
  wire  _T_1 = io_rd == 5'h0; // @[RegisterFile.scala 27:16]
  wire [31:0] _GEN_129 = 5'h1 == io_rd ? RegFile_1 : RegFile_0; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_130 = 5'h2 == io_rd ? RegFile_2 : _GEN_129; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_131 = 5'h3 == io_rd ? RegFile_3 : _GEN_130; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_132 = 5'h4 == io_rd ? RegFile_4 : _GEN_131; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_133 = 5'h5 == io_rd ? RegFile_5 : _GEN_132; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_134 = 5'h6 == io_rd ? RegFile_6 : _GEN_133; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_135 = 5'h7 == io_rd ? RegFile_7 : _GEN_134; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_136 = 5'h8 == io_rd ? RegFile_8 : _GEN_135; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_137 = 5'h9 == io_rd ? RegFile_9 : _GEN_136; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_138 = 5'ha == io_rd ? RegFile_10 : _GEN_137; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_139 = 5'hb == io_rd ? RegFile_11 : _GEN_138; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_140 = 5'hc == io_rd ? RegFile_12 : _GEN_139; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_141 = 5'hd == io_rd ? RegFile_13 : _GEN_140; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_142 = 5'he == io_rd ? RegFile_14 : _GEN_141; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_143 = 5'hf == io_rd ? RegFile_15 : _GEN_142; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_144 = 5'h10 == io_rd ? RegFile_16 : _GEN_143; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_145 = 5'h11 == io_rd ? RegFile_17 : _GEN_144; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_146 = 5'h12 == io_rd ? RegFile_18 : _GEN_145; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_147 = 5'h13 == io_rd ? RegFile_19 : _GEN_146; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_148 = 5'h14 == io_rd ? RegFile_20 : _GEN_147; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_149 = 5'h15 == io_rd ? RegFile_21 : _GEN_148; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_150 = 5'h16 == io_rd ? RegFile_22 : _GEN_149; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_151 = 5'h17 == io_rd ? RegFile_23 : _GEN_150; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_152 = 5'h18 == io_rd ? RegFile_24 : _GEN_151; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_153 = 5'h19 == io_rd ? RegFile_25 : _GEN_152; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_154 = 5'h1a == io_rd ? RegFile_26 : _GEN_153; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_155 = 5'h1b == io_rd ? RegFile_27 : _GEN_154; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_156 = 5'h1c == io_rd ? RegFile_28 : _GEN_155; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_157 = 5'h1d == io_rd ? RegFile_29 : _GEN_156; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_158 = 5'h1e == io_rd ? RegFile_30 : _GEN_157; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_159 = 5'h1f == io_rd ? RegFile_31 : _GEN_158; // @[RegisterFile.scala 31:{20,20}]
  wire [31:0] _GEN_96 = 5'h0 == io_rd ? _GEN_159 : RegFile_0; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_97 = 5'h1 == io_rd ? _GEN_159 : RegFile_1; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_98 = 5'h2 == io_rd ? _GEN_159 : RegFile_2; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_99 = 5'h3 == io_rd ? _GEN_159 : RegFile_3; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_100 = 5'h4 == io_rd ? _GEN_159 : RegFile_4; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_101 = 5'h5 == io_rd ? _GEN_159 : RegFile_5; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_102 = 5'h6 == io_rd ? _GEN_159 : RegFile_6; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_103 = 5'h7 == io_rd ? _GEN_159 : RegFile_7; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_104 = 5'h8 == io_rd ? _GEN_159 : RegFile_8; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_105 = 5'h9 == io_rd ? _GEN_159 : RegFile_9; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_106 = 5'ha == io_rd ? _GEN_159 : RegFile_10; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_107 = 5'hb == io_rd ? _GEN_159 : RegFile_11; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_108 = 5'hc == io_rd ? _GEN_159 : RegFile_12; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_109 = 5'hd == io_rd ? _GEN_159 : RegFile_13; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_110 = 5'he == io_rd ? _GEN_159 : RegFile_14; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_111 = 5'hf == io_rd ? _GEN_159 : RegFile_15; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_112 = 5'h10 == io_rd ? _GEN_159 : RegFile_16; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_113 = 5'h11 == io_rd ? _GEN_159 : RegFile_17; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_114 = 5'h12 == io_rd ? _GEN_159 : RegFile_18; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_115 = 5'h13 == io_rd ? _GEN_159 : RegFile_19; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_116 = 5'h14 == io_rd ? _GEN_159 : RegFile_20; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_117 = 5'h15 == io_rd ? _GEN_159 : RegFile_21; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_118 = 5'h16 == io_rd ? _GEN_159 : RegFile_22; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_119 = 5'h17 == io_rd ? _GEN_159 : RegFile_23; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_120 = 5'h18 == io_rd ? _GEN_159 : RegFile_24; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_121 = 5'h19 == io_rd ? _GEN_159 : RegFile_25; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_122 = 5'h1a == io_rd ? _GEN_159 : RegFile_26; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_123 = 5'h1b == io_rd ? _GEN_159 : RegFile_27; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_124 = 5'h1c == io_rd ? _GEN_159 : RegFile_28; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_125 = 5'h1d == io_rd ? _GEN_159 : RegFile_29; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_126 = 5'h1e == io_rd ? _GEN_159 : RegFile_30; // @[RegisterFile.scala 31:{20,20} 19:25]
  wire [31:0] _GEN_127 = 5'h1f == io_rd ? _GEN_159 : RegFile_31; // @[RegisterFile.scala 31:{20,20} 19:25]
  reg [31:0] io_operand1_REG; // @[RegisterFile.scala 37:25]
  wire [31:0] _GEN_257 = 5'h1 == io_rs1 ? RegFile_1 : RegFile_0; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_258 = 5'h2 == io_rs1 ? RegFile_2 : _GEN_257; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_259 = 5'h3 == io_rs1 ? RegFile_3 : _GEN_258; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_260 = 5'h4 == io_rs1 ? RegFile_4 : _GEN_259; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_261 = 5'h5 == io_rs1 ? RegFile_5 : _GEN_260; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_262 = 5'h6 == io_rs1 ? RegFile_6 : _GEN_261; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_263 = 5'h7 == io_rs1 ? RegFile_7 : _GEN_262; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_264 = 5'h8 == io_rs1 ? RegFile_8 : _GEN_263; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_265 = 5'h9 == io_rs1 ? RegFile_9 : _GEN_264; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_266 = 5'ha == io_rs1 ? RegFile_10 : _GEN_265; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_267 = 5'hb == io_rs1 ? RegFile_11 : _GEN_266; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_268 = 5'hc == io_rs1 ? RegFile_12 : _GEN_267; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_269 = 5'hd == io_rs1 ? RegFile_13 : _GEN_268; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_270 = 5'he == io_rs1 ? RegFile_14 : _GEN_269; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_271 = 5'hf == io_rs1 ? RegFile_15 : _GEN_270; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_272 = 5'h10 == io_rs1 ? RegFile_16 : _GEN_271; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_273 = 5'h11 == io_rs1 ? RegFile_17 : _GEN_272; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_274 = 5'h12 == io_rs1 ? RegFile_18 : _GEN_273; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_275 = 5'h13 == io_rs1 ? RegFile_19 : _GEN_274; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_276 = 5'h14 == io_rs1 ? RegFile_20 : _GEN_275; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_277 = 5'h15 == io_rs1 ? RegFile_21 : _GEN_276; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_278 = 5'h16 == io_rs1 ? RegFile_22 : _GEN_277; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_279 = 5'h17 == io_rs1 ? RegFile_23 : _GEN_278; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_280 = 5'h18 == io_rs1 ? RegFile_24 : _GEN_279; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_281 = 5'h19 == io_rs1 ? RegFile_25 : _GEN_280; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_282 = 5'h1a == io_rs1 ? RegFile_26 : _GEN_281; // @[RegisterFile.scala 37:{25,25}]
  wire [31:0] _GEN_283 = 5'h1b == io_rs1 ? RegFile_27 : _GEN_282; // @[RegisterFile.scala 37:{25,25}]
  reg [31:0] io_operand2_REG; // @[RegisterFile.scala 38:25]
  wire [31:0] _GEN_289 = 5'h1 == io_rs2 ? RegFile_1 : RegFile_0; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_290 = 5'h2 == io_rs2 ? RegFile_2 : _GEN_289; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_291 = 5'h3 == io_rs2 ? RegFile_3 : _GEN_290; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_292 = 5'h4 == io_rs2 ? RegFile_4 : _GEN_291; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_293 = 5'h5 == io_rs2 ? RegFile_5 : _GEN_292; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_294 = 5'h6 == io_rs2 ? RegFile_6 : _GEN_293; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_295 = 5'h7 == io_rs2 ? RegFile_7 : _GEN_294; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_296 = 5'h8 == io_rs2 ? RegFile_8 : _GEN_295; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_297 = 5'h9 == io_rs2 ? RegFile_9 : _GEN_296; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_298 = 5'ha == io_rs2 ? RegFile_10 : _GEN_297; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_299 = 5'hb == io_rs2 ? RegFile_11 : _GEN_298; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_300 = 5'hc == io_rs2 ? RegFile_12 : _GEN_299; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_301 = 5'hd == io_rs2 ? RegFile_13 : _GEN_300; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_302 = 5'he == io_rs2 ? RegFile_14 : _GEN_301; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_303 = 5'hf == io_rs2 ? RegFile_15 : _GEN_302; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_304 = 5'h10 == io_rs2 ? RegFile_16 : _GEN_303; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_305 = 5'h11 == io_rs2 ? RegFile_17 : _GEN_304; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_306 = 5'h12 == io_rs2 ? RegFile_18 : _GEN_305; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_307 = 5'h13 == io_rs2 ? RegFile_19 : _GEN_306; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_308 = 5'h14 == io_rs2 ? RegFile_20 : _GEN_307; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_309 = 5'h15 == io_rs2 ? RegFile_21 : _GEN_308; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_310 = 5'h16 == io_rs2 ? RegFile_22 : _GEN_309; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_311 = 5'h17 == io_rs2 ? RegFile_23 : _GEN_310; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_312 = 5'h18 == io_rs2 ? RegFile_24 : _GEN_311; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_313 = 5'h19 == io_rs2 ? RegFile_25 : _GEN_312; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_314 = 5'h1a == io_rs2 ? RegFile_26 : _GEN_313; // @[RegisterFile.scala 38:{25,25}]
  wire [31:0] _GEN_315 = 5'h1b == io_rs2 ? RegFile_27 : _GEN_314; // @[RegisterFile.scala 38:{25,25}]
  assign io_operand1 = io_operand1_REG; // @[RegisterFile.scala 37:15]
  assign io_operand2 = io_operand2_REG; // @[RegisterFile.scala 38:15]
  always @(posedge clock) begin
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_0 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h0 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_0 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_0 <= _GEN_0;
        end
      end else begin
        RegFile_0 <= _GEN_0;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h0 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_0 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_0 <= _GEN_96;
      end
    end else begin
      RegFile_0 <= _GEN_96;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_1 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_1 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_1 <= _GEN_1;
        end
      end else begin
        RegFile_1 <= _GEN_1;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_1 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_1 <= _GEN_97;
      end
    end else begin
      RegFile_1 <= _GEN_97;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_2 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h2 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_2 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_2 <= _GEN_2;
        end
      end else begin
        RegFile_2 <= _GEN_2;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h2 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_2 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_2 <= _GEN_98;
      end
    end else begin
      RegFile_2 <= _GEN_98;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_3 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h3 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_3 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_3 <= _GEN_3;
        end
      end else begin
        RegFile_3 <= _GEN_3;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h3 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_3 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_3 <= _GEN_99;
      end
    end else begin
      RegFile_3 <= _GEN_99;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_4 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h4 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_4 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_4 <= _GEN_4;
        end
      end else begin
        RegFile_4 <= _GEN_4;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h4 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_4 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_4 <= _GEN_100;
      end
    end else begin
      RegFile_4 <= _GEN_100;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_5 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h5 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_5 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_5 <= _GEN_5;
        end
      end else begin
        RegFile_5 <= _GEN_5;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h5 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_5 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_5 <= _GEN_101;
      end
    end else begin
      RegFile_5 <= _GEN_101;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_6 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h6 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_6 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_6 <= _GEN_6;
        end
      end else begin
        RegFile_6 <= _GEN_6;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h6 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_6 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_6 <= _GEN_102;
      end
    end else begin
      RegFile_6 <= _GEN_102;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_7 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h7 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_7 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_7 <= _GEN_7;
        end
      end else begin
        RegFile_7 <= _GEN_7;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h7 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_7 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_7 <= _GEN_103;
      end
    end else begin
      RegFile_7 <= _GEN_103;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_8 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h8 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_8 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_8 <= _GEN_8;
        end
      end else begin
        RegFile_8 <= _GEN_8;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h8 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_8 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_8 <= _GEN_104;
      end
    end else begin
      RegFile_8 <= _GEN_104;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_9 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h9 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_9 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_9 <= _GEN_9;
        end
      end else begin
        RegFile_9 <= _GEN_9;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h9 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_9 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_9 <= _GEN_105;
      end
    end else begin
      RegFile_9 <= _GEN_105;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_10 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'ha == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_10 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_10 <= _GEN_10;
        end
      end else begin
        RegFile_10 <= _GEN_10;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'ha == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_10 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_10 <= _GEN_106;
      end
    end else begin
      RegFile_10 <= _GEN_106;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_11 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'hb == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_11 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_11 <= _GEN_11;
        end
      end else begin
        RegFile_11 <= _GEN_11;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'hb == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_11 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_11 <= _GEN_107;
      end
    end else begin
      RegFile_11 <= _GEN_107;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_12 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'hc == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_12 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_12 <= _GEN_12;
        end
      end else begin
        RegFile_12 <= _GEN_12;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'hc == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_12 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_12 <= _GEN_108;
      end
    end else begin
      RegFile_12 <= _GEN_108;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_13 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'hd == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_13 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_13 <= _GEN_13;
        end
      end else begin
        RegFile_13 <= _GEN_13;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'hd == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_13 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_13 <= _GEN_109;
      end
    end else begin
      RegFile_13 <= _GEN_109;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_14 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'he == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_14 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_14 <= _GEN_14;
        end
      end else begin
        RegFile_14 <= _GEN_14;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'he == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_14 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_14 <= _GEN_110;
      end
    end else begin
      RegFile_14 <= _GEN_110;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_15 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'hf == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_15 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_15 <= _GEN_15;
        end
      end else begin
        RegFile_15 <= _GEN_15;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'hf == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_15 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_15 <= _GEN_111;
      end
    end else begin
      RegFile_15 <= _GEN_111;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_16 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h10 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_16 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_16 <= _GEN_16;
        end
      end else begin
        RegFile_16 <= _GEN_16;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h10 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_16 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_16 <= _GEN_112;
      end
    end else begin
      RegFile_16 <= _GEN_112;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_17 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h11 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_17 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_17 <= _GEN_17;
        end
      end else begin
        RegFile_17 <= _GEN_17;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h11 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_17 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_17 <= _GEN_113;
      end
    end else begin
      RegFile_17 <= _GEN_113;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_18 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h12 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_18 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_18 <= _GEN_18;
        end
      end else begin
        RegFile_18 <= _GEN_18;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h12 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_18 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_18 <= _GEN_114;
      end
    end else begin
      RegFile_18 <= _GEN_114;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_19 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h13 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_19 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_19 <= _GEN_19;
        end
      end else begin
        RegFile_19 <= _GEN_19;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h13 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_19 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_19 <= _GEN_115;
      end
    end else begin
      RegFile_19 <= _GEN_115;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_20 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h14 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_20 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_20 <= _GEN_20;
        end
      end else begin
        RegFile_20 <= _GEN_20;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h14 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_20 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_20 <= _GEN_116;
      end
    end else begin
      RegFile_20 <= _GEN_116;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_21 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h15 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_21 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_21 <= _GEN_21;
        end
      end else begin
        RegFile_21 <= _GEN_21;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h15 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_21 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_21 <= _GEN_117;
      end
    end else begin
      RegFile_21 <= _GEN_117;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_22 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h16 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_22 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_22 <= _GEN_22;
        end
      end else begin
        RegFile_22 <= _GEN_22;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h16 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_22 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_22 <= _GEN_118;
      end
    end else begin
      RegFile_22 <= _GEN_118;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_23 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h17 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_23 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_23 <= _GEN_23;
        end
      end else begin
        RegFile_23 <= _GEN_23;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h17 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_23 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_23 <= _GEN_119;
      end
    end else begin
      RegFile_23 <= _GEN_119;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_24 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h18 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_24 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_24 <= _GEN_24;
        end
      end else begin
        RegFile_24 <= _GEN_24;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h18 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_24 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_24 <= _GEN_120;
      end
    end else begin
      RegFile_24 <= _GEN_120;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_25 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h19 == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_25 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_25 <= _GEN_25;
        end
      end else begin
        RegFile_25 <= _GEN_25;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h19 == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_25 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_25 <= _GEN_121;
      end
    end else begin
      RegFile_25 <= _GEN_121;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_26 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1a == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_26 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_26 <= _GEN_26;
        end
      end else begin
        RegFile_26 <= _GEN_26;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1a == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_26 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_26 <= _GEN_122;
      end
    end else begin
      RegFile_26 <= _GEN_122;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_27 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1b == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_27 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_27 <= _GEN_27;
        end
      end else begin
        RegFile_27 <= _GEN_27;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1b == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_27 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_27 <= _GEN_123;
      end
    end else begin
      RegFile_27 <= _GEN_123;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_28 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1c == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_28 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_28 <= _GEN_28;
        end
      end else begin
        RegFile_28 <= _GEN_28;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1c == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_28 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_28 <= _GEN_124;
      end
    end else begin
      RegFile_28 <= _GEN_124;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_29 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1d == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_29 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_29 <= _GEN_29;
        end
      end else begin
        RegFile_29 <= _GEN_29;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1d == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_29 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_29 <= _GEN_125;
      end
    end else begin
      RegFile_29 <= _GEN_125;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_30 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1e == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_30 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_30 <= _GEN_30;
        end
      end else begin
        RegFile_30 <= _GEN_30;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1e == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_30 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_30 <= _GEN_126;
      end
    end else begin
      RegFile_30 <= _GEN_126;
    end
    if (reset) begin // @[RegisterFile.scala 19:25]
      RegFile_31 <= 32'h0; // @[RegisterFile.scala 19:25]
    end else if (io_writeEnable) begin // @[RegisterFile.scala 25:33]
      if (io_rd == 5'h0) begin // @[RegisterFile.scala 27:24]
        if (5'h1f == io_rd) begin // @[RegisterFile.scala 28:22]
          RegFile_31 <= 32'h0; // @[RegisterFile.scala 28:22]
        end else begin
          RegFile_31 <= _GEN_31;
        end
      end else begin
        RegFile_31 <= _GEN_31;
      end
    end else if (_T_1) begin // @[RegisterFile.scala 32:25]
      if (5'h1f == io_rd) begin // @[RegisterFile.scala 33:22]
        RegFile_31 <= 32'h0; // @[RegisterFile.scala 33:22]
      end else begin
        RegFile_31 <= _GEN_127;
      end
    end else begin
      RegFile_31 <= _GEN_127;
    end
    if (5'h1f == io_rs1) begin // @[RegisterFile.scala 37:25]
      io_operand1_REG <= RegFile_31; // @[RegisterFile.scala 37:25]
    end else if (5'h1e == io_rs1) begin // @[RegisterFile.scala 37:25]
      io_operand1_REG <= RegFile_30; // @[RegisterFile.scala 37:25]
    end else if (5'h1d == io_rs1) begin // @[RegisterFile.scala 37:25]
      io_operand1_REG <= RegFile_29; // @[RegisterFile.scala 37:25]
    end else if (5'h1c == io_rs1) begin // @[RegisterFile.scala 37:25]
      io_operand1_REG <= RegFile_28; // @[RegisterFile.scala 37:25]
    end else begin
      io_operand1_REG <= _GEN_283;
    end
    if (5'h1f == io_rs2) begin // @[RegisterFile.scala 38:25]
      io_operand2_REG <= RegFile_31; // @[RegisterFile.scala 38:25]
    end else if (5'h1e == io_rs2) begin // @[RegisterFile.scala 38:25]
      io_operand2_REG <= RegFile_30; // @[RegisterFile.scala 38:25]
    end else if (5'h1d == io_rs2) begin // @[RegisterFile.scala 38:25]
      io_operand2_REG <= RegFile_29; // @[RegisterFile.scala 38:25]
    end else if (5'h1c == io_rs2) begin // @[RegisterFile.scala 38:25]
      io_operand2_REG <= RegFile_28; // @[RegisterFile.scala 38:25]
    end else begin
      io_operand2_REG <= _GEN_315;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegFile_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  RegFile_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  RegFile_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  RegFile_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  RegFile_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  RegFile_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  RegFile_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  RegFile_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  RegFile_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  RegFile_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  RegFile_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  RegFile_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  RegFile_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  RegFile_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  RegFile_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  RegFile_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  RegFile_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  RegFile_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  RegFile_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  RegFile_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  RegFile_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  RegFile_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  RegFile_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  RegFile_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  RegFile_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  RegFile_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  RegFile_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  RegFile_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  RegFile_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  RegFile_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  RegFile_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  RegFile_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  io_operand1_REG = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  io_operand2_REG = _RAND_33[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ImmediateGenerator(
  input  [2:0]  io_instrType,
  input  [31:0] io_instruction,
  output [31:0] io_immediate
);
  wire [19:0] _io_immediate_T_2 = io_instruction[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _io_immediate_T_4 = {_io_immediate_T_2,io_instruction[31:20]}; // @[Cat.scala 33:92]
  wire [11:0] _io_immediate_T_7 = {io_instruction[31:25],io_instruction[11:7]}; // @[Cat.scala 33:92]
  wire [12:0] _io_immediate_T_12 = {io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8],1'h0
    }; // @[Cat.scala 33:92]
  wire [31:0] _io_immediate_T_14 = {io_instruction[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [20:0] _io_immediate_T_19 = {io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:21],1'h0
    }; // @[Cat.scala 33:92]
  wire [31:0] _GEN_0 = 3'h5 == io_instrType ? {{11'd0}, _io_immediate_T_19} : 32'h0; // @[ImmediateGenerator.scala 13:16 14:23 31:20]
  wire [31:0] _GEN_1 = 3'h4 == io_instrType ? _io_immediate_T_14 : _GEN_0; // @[ImmediateGenerator.scala 14:23 28:20]
  wire [31:0] _GEN_2 = 3'h3 == io_instrType ? {{19'd0}, _io_immediate_T_12} : _GEN_1; // @[ImmediateGenerator.scala 14:23 25:20]
  wire [31:0] _GEN_3 = 3'h2 == io_instrType ? {{20'd0}, _io_immediate_T_7} : _GEN_2; // @[ImmediateGenerator.scala 14:23 22:20]
  wire [31:0] _GEN_4 = 3'h1 == io_instrType ? _io_immediate_T_4 : _GEN_3; // @[ImmediateGenerator.scala 14:23 19:20]
  assign io_immediate = 3'h0 == io_instrType ? 32'h0 : _GEN_4; // @[ImmediateGenerator.scala 14:23 16:20]
endmodule
module ControlUnit(
  input  [2:0] io_funct3,
  input  [6:0] io_funct7,
  input  [6:0] io_opcode,
  output       io_MuxAluSel,
  output [7:0] io_AluSel,
  output       io_RegWriteEnable,
  output       io_WriteDataMux,
  output       io_MemWriteEnable
);
  wire [9:0] io_AluSel_compositeKey = {io_funct3,io_funct7}; // @[Cat.scala 33:92]
  wire [2:0] _io_AluSel_T_15 = 10'h200 == io_AluSel_compositeKey ? 3'h4 : {{2'd0}, 10'h20 == io_AluSel_compositeKey}; // @[Mux.scala 81:58]
  wire [2:0] _io_AluSel_T_17 = 10'h300 == io_AluSel_compositeKey ? 3'h3 : _io_AluSel_T_15; // @[Mux.scala 81:58]
  wire [2:0] _io_AluSel_T_19 = 10'h380 == io_AluSel_compositeKey ? 3'h2 : _io_AluSel_T_17; // @[Mux.scala 81:58]
  wire [2:0] _io_AluSel_T_21 = 10'h80 == io_AluSel_compositeKey ? 3'h5 : _io_AluSel_T_19; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_23 = 10'h100 == io_AluSel_compositeKey ? 4'h8 : {{1'd0}, _io_AluSel_T_21}; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_25 = 10'h180 == io_AluSel_compositeKey ? 4'h9 : _io_AluSel_T_23; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_27 = 10'h280 == io_AluSel_compositeKey ? 4'h6 : _io_AluSel_T_25; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_29 = 10'h2a0 == io_AluSel_compositeKey ? 4'h7 : _io_AluSel_T_27; // @[Mux.scala 81:58]
  wire  _io_MuxAluSel_T_1 = io_opcode == 7'h33 ? 1'h0 : 1'h1; // @[ControlUnit.scala 54:26]
  wire [3:0] _io_AluSel_T_31 = 3'h0 == io_funct3 ? 4'ha : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_33 = 3'h1 == io_funct3 ? 4'hb : _io_AluSel_T_31; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_35 = 3'h4 == io_funct3 ? 4'hc : _io_AluSel_T_33; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_37 = 3'h5 == io_funct3 ? 4'hd : _io_AluSel_T_35; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_39 = 3'h6 == io_funct3 ? 4'he : _io_AluSel_T_37; // @[Mux.scala 81:58]
  wire [3:0] _io_AluSel_T_41 = 3'h7 == io_funct3 ? 4'hf : _io_AluSel_T_39; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_43 = 3'h0 == io_funct3 ? 5'h10 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_45 = 3'h1 == io_funct3 ? 5'h11 : _io_AluSel_T_43; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_47 = 3'h2 == io_funct3 ? 5'h12 : _io_AluSel_T_45; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_49 = 3'h4 == io_funct3 ? 5'h13 : _io_AluSel_T_47; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_51 = 3'h5 == io_funct3 ? 5'h14 : _io_AluSel_T_49; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_53 = 3'h0 == io_funct3 ? 5'h15 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_55 = 3'h1 == io_funct3 ? 5'h16 : _io_AluSel_T_53; // @[Mux.scala 81:58]
  wire [4:0] _io_AluSel_T_57 = 3'h2 == io_funct3 ? 5'h17 : _io_AluSel_T_55; // @[Mux.scala 81:58]
  wire [4:0] _GEN_2 = 7'h23 == io_opcode ? _io_AluSel_T_57 : 5'h0; // @[ControlUnit.scala 27:13 50:21 84:17]
  wire [4:0] _GEN_5 = 7'h3 == io_opcode ? _io_AluSel_T_51 : _GEN_2; // @[ControlUnit.scala 50:21 72:17]
  wire  _GEN_6 = 7'h3 == io_opcode ? 1'h0 : 7'h23 == io_opcode; // @[ControlUnit.scala 23:21 50:21]
  wire  _GEN_7 = 7'h63 == io_opcode ? 1'h0 : 7'h3 == io_opcode; // @[ControlUnit.scala 50:21 58:25]
  wire [4:0] _GEN_8 = 7'h63 == io_opcode ? {{1'd0}, _io_AluSel_T_41} : _GEN_5; // @[ControlUnit.scala 50:21 59:17]
  wire  _GEN_10 = 7'h63 == io_opcode ? 1'h0 : _GEN_6; // @[ControlUnit.scala 23:21 50:21]
  wire [4:0] _GEN_12 = 7'h33 == io_opcode | 7'h13 == io_opcode ? {{1'd0}, _io_AluSel_T_29} : _GEN_8; // @[ControlUnit.scala 50:21 53:17]
  assign io_MuxAluSel = 7'h33 == io_opcode | 7'h13 == io_opcode ? _io_MuxAluSel_T_1 : 1'h1; // @[ControlUnit.scala 28:16 50:21 54:20]
  assign io_AluSel = {{3'd0}, _GEN_12};
  assign io_RegWriteEnable = 7'h33 == io_opcode | 7'h13 == io_opcode | _GEN_7; // @[ControlUnit.scala 50:21 52:25]
  assign io_WriteDataMux = 7'h33 == io_opcode | 7'h13 == io_opcode ? 1'h0 : _GEN_7; // @[ControlUnit.scala 26:19 50:21]
  assign io_MemWriteEnable = 7'h33 == io_opcode | 7'h13 == io_opcode ? 1'h0 : _GEN_10; // @[ControlUnit.scala 23:21 50:21]
endmodule
module ALU(
  input  [7:0]  io_ALUSel,
  input  [31:0] io_operand1,
  input  [31:0] io_operand2,
  output [31:0] io_ALURes
);
  wire [31:0] signedOperand2 = io_operand2; // @[ALU.scala 17:36]
  wire [31:0] _io_ALURes_T_3 = $signed(io_operand1) + $signed(io_operand2); // @[ALU.scala 23:54]
  wire [31:0] _io_ALURes_T_7 = $signed(io_operand1) - $signed(io_operand2); // @[ALU.scala 26:54]
  wire [31:0] _io_ALURes_T_10 = $signed(io_operand1) & $signed(io_operand2); // @[ALU.scala 29:54]
  wire [31:0] _io_ALURes_T_13 = $signed(io_operand1) | $signed(io_operand2); // @[ALU.scala 32:54]
  wire [31:0] _io_ALURes_T_16 = $signed(io_operand1) ^ $signed(io_operand2); // @[ALU.scala 35:54]
  wire [62:0] _GEN_0 = {{31'd0}, io_operand1}; // @[ALU.scala 38:33]
  wire [62:0] _io_ALURes_T_18 = _GEN_0 << io_operand2[4:0]; // @[ALU.scala 38:33]
  wire [31:0] _io_ALURes_T_20 = io_operand1 >> io_operand2[4:0]; // @[ALU.scala 41:33]
  wire [31:0] _io_ALURes_T_23 = $signed(io_operand1) >>> signedOperand2[4:0]; // @[ALU.scala 45:62]
  wire  _T_9 = $signed(io_operand1) < $signed(io_operand2); // @[ALU.scala 48:27]
  wire  _T_11 = io_operand1 < io_operand2; // @[ALU.scala 55:24]
  wire [5:0] _GEN_2 = 8'h9 == io_ALUSel ? {{5'd0}, _T_11} : 6'h2a; // @[ALU.scala 20:13 21:21]
  wire [5:0] _GEN_3 = 8'h8 == io_ALUSel ? {{5'd0}, _T_9} : _GEN_2; // @[ALU.scala 21:21]
  wire [31:0] _GEN_4 = 8'h7 == io_ALUSel ? _io_ALURes_T_23 : {{26'd0}, _GEN_3}; // @[ALU.scala 21:21 45:17]
  wire [31:0] _GEN_5 = 8'h6 == io_ALUSel ? _io_ALURes_T_20 : _GEN_4; // @[ALU.scala 21:21 41:17]
  wire [62:0] _GEN_6 = 8'h5 == io_ALUSel ? _io_ALURes_T_18 : {{31'd0}, _GEN_5}; // @[ALU.scala 21:21 38:17]
  wire [62:0] _GEN_7 = 8'h4 == io_ALUSel ? {{31'd0}, _io_ALURes_T_16} : _GEN_6; // @[ALU.scala 21:21 35:17]
  wire [62:0] _GEN_8 = 8'h3 == io_ALUSel ? {{31'd0}, _io_ALURes_T_13} : _GEN_7; // @[ALU.scala 21:21 32:17]
  wire [62:0] _GEN_9 = 8'h2 == io_ALUSel ? {{31'd0}, _io_ALURes_T_10} : _GEN_8; // @[ALU.scala 21:21 29:17]
  wire [62:0] _GEN_10 = 8'h1 == io_ALUSel ? {{31'd0}, _io_ALURes_T_7} : _GEN_9; // @[ALU.scala 21:21 26:17]
  wire [62:0] _GEN_11 = 8'h0 == io_ALUSel ? {{31'd0}, _io_ALURes_T_3} : _GEN_10; // @[ALU.scala 21:21 23:17]
  assign io_ALURes = _GEN_11[31:0];
endmodule
module EXStage(
  input         clock,
  input         reset,
  input  [31:0] io_instruction,
  input  [2:0]  io_instrType,
  input  [2:0]  io_funct3,
  input  [6:0]  io_funct7,
  input  [6:0]  io_opcode,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [31:0] io_writeData,
  input         io_writeEnable,
  input  [4:0]  io_rdReg,
  output [31:0] io_ALURes,
  output [31:0] io_address,
  output [31:0] io_dataWriteMem,
  output [4:0]  io_rdRegIn,
  output        io_RegWriteEnable,
  output        io_WriteDataMux,
  output        io_MemWriteEnable,
  output        io_readIsIO,
  output        io_IOWriteEnable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  RegFile_clock; // @[EXStage.scala 34:23]
  wire  RegFile_reset; // @[EXStage.scala 34:23]
  wire [4:0] RegFile_io_rs1; // @[EXStage.scala 34:23]
  wire [4:0] RegFile_io_rs2; // @[EXStage.scala 34:23]
  wire [31:0] RegFile_io_writeData; // @[EXStage.scala 34:23]
  wire [4:0] RegFile_io_rd; // @[EXStage.scala 34:23]
  wire  RegFile_io_writeEnable; // @[EXStage.scala 34:23]
  wire [31:0] RegFile_io_operand1; // @[EXStage.scala 34:23]
  wire [31:0] RegFile_io_operand2; // @[EXStage.scala 34:23]
  wire [2:0] immGen_io_instrType; // @[EXStage.scala 35:22]
  wire [31:0] immGen_io_instruction; // @[EXStage.scala 35:22]
  wire [31:0] immGen_io_immediate; // @[EXStage.scala 35:22]
  wire [2:0] controlUnit_io_funct3; // @[EXStage.scala 36:27]
  wire [6:0] controlUnit_io_funct7; // @[EXStage.scala 36:27]
  wire [6:0] controlUnit_io_opcode; // @[EXStage.scala 36:27]
  wire  controlUnit_io_MuxAluSel; // @[EXStage.scala 36:27]
  wire [7:0] controlUnit_io_AluSel; // @[EXStage.scala 36:27]
  wire  controlUnit_io_RegWriteEnable; // @[EXStage.scala 36:27]
  wire  controlUnit_io_WriteDataMux; // @[EXStage.scala 36:27]
  wire  controlUnit_io_MemWriteEnable; // @[EXStage.scala 36:27]
  wire [7:0] ALU_io_ALUSel; // @[EXStage.scala 37:19]
  wire [31:0] ALU_io_operand1; // @[EXStage.scala 37:19]
  wire [31:0] ALU_io_operand2; // @[EXStage.scala 37:19]
  wire [31:0] ALU_io_ALURes; // @[EXStage.scala 37:19]
  reg [31:0] instructionReg; // @[EXStage.scala 40:31]
  reg [2:0] instrTypeReg; // @[EXStage.scala 41:29]
  reg [2:0] funct3Reg; // @[EXStage.scala 42:26]
  reg [6:0] funct7Reg; // @[EXStage.scala 43:26]
  reg [6:0] opcodeReg; // @[EXStage.scala 44:26]
  reg [4:0] rdReg; // @[EXStage.scala 45:22]
  RegisterFile RegFile ( // @[EXStage.scala 34:23]
    .clock(RegFile_clock),
    .reset(RegFile_reset),
    .io_rs1(RegFile_io_rs1),
    .io_rs2(RegFile_io_rs2),
    .io_writeData(RegFile_io_writeData),
    .io_rd(RegFile_io_rd),
    .io_writeEnable(RegFile_io_writeEnable),
    .io_operand1(RegFile_io_operand1),
    .io_operand2(RegFile_io_operand2)
  );
  ImmediateGenerator immGen ( // @[EXStage.scala 35:22]
    .io_instrType(immGen_io_instrType),
    .io_instruction(immGen_io_instruction),
    .io_immediate(immGen_io_immediate)
  );
  ControlUnit controlUnit ( // @[EXStage.scala 36:27]
    .io_funct3(controlUnit_io_funct3),
    .io_funct7(controlUnit_io_funct7),
    .io_opcode(controlUnit_io_opcode),
    .io_MuxAluSel(controlUnit_io_MuxAluSel),
    .io_AluSel(controlUnit_io_AluSel),
    .io_RegWriteEnable(controlUnit_io_RegWriteEnable),
    .io_WriteDataMux(controlUnit_io_WriteDataMux),
    .io_MemWriteEnable(controlUnit_io_MemWriteEnable)
  );
  ALU ALU ( // @[EXStage.scala 37:19]
    .io_ALUSel(ALU_io_ALUSel),
    .io_operand1(ALU_io_operand1),
    .io_operand2(ALU_io_operand2),
    .io_ALURes(ALU_io_ALURes)
  );
  assign io_ALURes = ALU_io_ALURes; // @[EXStage.scala 80:15]
  assign io_address = ALU_io_ALURes; // @[EXStage.scala 81:14]
  assign io_dataWriteMem = RegFile_io_operand2; // @[EXStage.scala 75:19]
  assign io_rdRegIn = rdReg; // @[EXStage.scala 110:14]
  assign io_RegWriteEnable = controlUnit_io_RegWriteEnable; // @[EXStage.scala 94:21]
  assign io_WriteDataMux = controlUnit_io_WriteDataMux; // @[EXStage.scala 95:19]
  assign io_MemWriteEnable = ALU_io_ALURes >= 32'h400 ? 1'h0 : controlUnit_io_MemWriteEnable; // @[EXStage.scala 102:33 103:23 97:21]
  assign io_readIsIO = ALU_io_ALURes >= 32'h400; // @[EXStage.scala 102:22]
  assign io_IOWriteEnable = ALU_io_ALURes >= 32'h400 & controlUnit_io_MemWriteEnable; // @[EXStage.scala 102:33 105:22 67:20]
  assign RegFile_clock = clock;
  assign RegFile_reset = reset;
  assign RegFile_io_rs1 = io_rs1; // @[EXStage.scala 70:18]
  assign RegFile_io_rs2 = io_rs2; // @[EXStage.scala 71:18]
  assign RegFile_io_writeData = io_writeData; // @[EXStage.scala 73:24]
  assign RegFile_io_rd = io_rdReg; // @[EXStage.scala 72:17]
  assign RegFile_io_writeEnable = io_writeEnable; // @[EXStage.scala 74:26]
  assign immGen_io_instrType = instrTypeReg; // @[EXStage.scala 84:23]
  assign immGen_io_instruction = instructionReg; // @[EXStage.scala 85:25]
  assign controlUnit_io_funct3 = funct3Reg; // @[EXStage.scala 89:25]
  assign controlUnit_io_funct7 = funct7Reg; // @[EXStage.scala 90:25]
  assign controlUnit_io_opcode = opcodeReg; // @[EXStage.scala 92:25]
  assign ALU_io_ALUSel = controlUnit_io_AluSel; // @[EXStage.scala 98:17]
  assign ALU_io_operand1 = RegFile_io_operand1; // @[EXStage.scala 78:19]
  assign ALU_io_operand2 = controlUnit_io_MuxAluSel ? immGen_io_immediate : RegFile_io_operand2; // @[EXStage.scala 79:25]
  always @(posedge clock) begin
    if (reset) begin // @[EXStage.scala 40:31]
      instructionReg <= 32'h0; // @[EXStage.scala 40:31]
    end else begin
      instructionReg <= io_instruction; // @[EXStage.scala 49:18]
    end
    if (reset) begin // @[EXStage.scala 41:29]
      instrTypeReg <= 3'h0; // @[EXStage.scala 41:29]
    end else begin
      instrTypeReg <= io_instrType; // @[EXStage.scala 50:16]
    end
    if (reset) begin // @[EXStage.scala 42:26]
      funct3Reg <= 3'h0; // @[EXStage.scala 42:26]
    end else begin
      funct3Reg <= io_funct3; // @[EXStage.scala 51:13]
    end
    if (reset) begin // @[EXStage.scala 43:26]
      funct7Reg <= 7'h0; // @[EXStage.scala 43:26]
    end else begin
      funct7Reg <= io_funct7; // @[EXStage.scala 52:13]
    end
    if (reset) begin // @[EXStage.scala 44:26]
      opcodeReg <= 7'h0; // @[EXStage.scala 44:26]
    end else begin
      opcodeReg <= io_opcode; // @[EXStage.scala 53:13]
    end
    if (reset) begin // @[EXStage.scala 45:22]
      rdReg <= 5'h0; // @[EXStage.scala 45:22]
    end else begin
      rdReg <= io_rd; // @[EXStage.scala 54:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instructionReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  instrTypeReg = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  funct3Reg = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  funct7Reg = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  opcodeReg = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  rdReg = _RAND_5[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataMemoryTest(
  input         clock,
  input         reset,
  input  [9:0]  io_addr,
  input         io_enableWrite,
  input  [31:0] io_dataIn,
  output [31:0] io_dataOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_2; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_3; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_4; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_5; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_6; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_7; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_8; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_9; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_10; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_11; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_12; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_13; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_14; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_15; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_16; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_17; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_18; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_19; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_20; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_21; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_22; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_23; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_24; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_25; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_26; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_27; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_28; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_29; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_30; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_31; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_32; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_33; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_34; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_35; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_36; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_37; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_38; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_39; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_40; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_41; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_42; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_43; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_44; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_45; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_46; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_47; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_48; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_49; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_50; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_51; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_52; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_53; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_54; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_55; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_56; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_57; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_58; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_59; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_60; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_61; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_62; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_63; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_64; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_65; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_66; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_67; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_68; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_69; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_70; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_71; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_72; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_73; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_74; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_75; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_76; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_77; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_78; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_79; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_80; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_81; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_82; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_83; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_84; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_85; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_86; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_87; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_88; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_89; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_90; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_91; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_92; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_93; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_94; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_95; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_96; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_97; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_98; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_99; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_100; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_101; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_102; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_103; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_104; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_105; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_106; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_107; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_108; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_109; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_110; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_111; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_112; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_113; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_114; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_115; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_116; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_117; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_118; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_119; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_120; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_121; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_122; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_123; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_124; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_125; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_126; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_127; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_128; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_129; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_130; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_131; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_132; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_133; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_134; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_135; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_136; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_137; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_138; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_139; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_140; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_141; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_142; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_143; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_144; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_145; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_146; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_147; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_148; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_149; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_150; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_151; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_152; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_153; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_154; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_155; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_156; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_157; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_158; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_159; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_160; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_161; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_162; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_163; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_164; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_165; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_166; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_167; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_168; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_169; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_170; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_171; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_172; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_173; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_174; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_175; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_176; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_177; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_178; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_179; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_180; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_181; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_182; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_183; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_184; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_185; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_186; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_187; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_188; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_189; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_190; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_191; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_192; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_193; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_194; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_195; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_196; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_197; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_198; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_199; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_200; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_201; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_202; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_203; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_204; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_205; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_206; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_207; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_208; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_209; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_210; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_211; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_212; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_213; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_214; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_215; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_216; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_217; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_218; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_219; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_220; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_221; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_222; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_223; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_224; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_225; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_226; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_227; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_228; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_229; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_230; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_231; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_232; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_233; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_234; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_235; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_236; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_237; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_238; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_239; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_240; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_241; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_242; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_243; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_244; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_245; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_246; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_247; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_248; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_249; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_250; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_251; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_252; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_253; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_254; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_255; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_256; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_257; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_258; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_259; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_260; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_261; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_262; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_263; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_264; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_265; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_266; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_267; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_268; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_269; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_270; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_271; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_272; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_273; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_274; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_275; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_276; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_277; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_278; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_279; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_280; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_281; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_282; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_283; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_284; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_285; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_286; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_287; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_288; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_289; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_290; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_291; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_292; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_293; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_294; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_295; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_296; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_297; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_298; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_299; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_300; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_301; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_302; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_303; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_304; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_305; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_306; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_307; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_308; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_309; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_310; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_311; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_312; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_313; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_314; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_315; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_316; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_317; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_318; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_319; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_320; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_321; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_322; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_323; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_324; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_325; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_326; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_327; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_328; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_329; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_330; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_331; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_332; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_333; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_334; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_335; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_336; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_337; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_338; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_339; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_340; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_341; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_342; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_343; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_344; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_345; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_346; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_347; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_348; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_349; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_350; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_351; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_352; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_353; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_354; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_355; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_356; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_357; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_358; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_359; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_360; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_361; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_362; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_363; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_364; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_365; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_366; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_367; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_368; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_369; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_370; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_371; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_372; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_373; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_374; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_375; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_376; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_377; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_378; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_379; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_380; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_381; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_382; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_383; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_384; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_385; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_386; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_387; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_388; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_389; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_390; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_391; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_392; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_393; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_394; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_395; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_396; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_397; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_398; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_399; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_400; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_401; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_402; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_403; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_404; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_405; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_406; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_407; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_408; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_409; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_410; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_411; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_412; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_413; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_414; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_415; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_416; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_417; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_418; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_419; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_420; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_421; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_422; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_423; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_424; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_425; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_426; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_427; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_428; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_429; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_430; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_431; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_432; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_433; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_434; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_435; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_436; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_437; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_438; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_439; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_440; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_441; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_442; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_443; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_444; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_445; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_446; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_447; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_448; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_449; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_450; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_451; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_452; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_453; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_454; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_455; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_456; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_457; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_458; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_459; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_460; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_461; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_462; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_463; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_464; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_465; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_466; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_467; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_468; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_469; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_470; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_471; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_472; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_473; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_474; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_475; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_476; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_477; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_478; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_479; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_480; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_481; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_482; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_483; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_484; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_485; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_486; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_487; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_488; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_489; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_490; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_491; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_492; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_493; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_494; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_495; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_496; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_497; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_498; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_499; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_500; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_501; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_502; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_503; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_504; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_505; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_506; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_507; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_508; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_509; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_510; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_511; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_512; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_513; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_514; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_515; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_516; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_517; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_518; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_519; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_520; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_521; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_522; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_523; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_524; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_525; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_526; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_527; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_528; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_529; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_530; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_531; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_532; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_533; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_534; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_535; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_536; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_537; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_538; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_539; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_540; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_541; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_542; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_543; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_544; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_545; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_546; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_547; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_548; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_549; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_550; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_551; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_552; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_553; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_554; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_555; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_556; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_557; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_558; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_559; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_560; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_561; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_562; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_563; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_564; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_565; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_566; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_567; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_568; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_569; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_570; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_571; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_572; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_573; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_574; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_575; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_576; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_577; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_578; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_579; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_580; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_581; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_582; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_583; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_584; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_585; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_586; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_587; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_588; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_589; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_590; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_591; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_592; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_593; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_594; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_595; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_596; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_597; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_598; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_599; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_600; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_601; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_602; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_603; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_604; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_605; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_606; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_607; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_608; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_609; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_610; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_611; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_612; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_613; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_614; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_615; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_616; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_617; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_618; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_619; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_620; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_621; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_622; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_623; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_624; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_625; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_626; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_627; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_628; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_629; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_630; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_631; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_632; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_633; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_634; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_635; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_636; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_637; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_638; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_639; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_640; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_641; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_642; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_643; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_644; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_645; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_646; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_647; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_648; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_649; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_650; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_651; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_652; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_653; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_654; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_655; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_656; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_657; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_658; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_659; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_660; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_661; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_662; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_663; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_664; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_665; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_666; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_667; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_668; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_669; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_670; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_671; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_672; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_673; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_674; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_675; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_676; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_677; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_678; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_679; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_680; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_681; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_682; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_683; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_684; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_685; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_686; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_687; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_688; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_689; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_690; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_691; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_692; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_693; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_694; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_695; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_696; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_697; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_698; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_699; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_700; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_701; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_702; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_703; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_704; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_705; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_706; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_707; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_708; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_709; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_710; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_711; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_712; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_713; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_714; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_715; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_716; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_717; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_718; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_719; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_720; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_721; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_722; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_723; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_724; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_725; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_726; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_727; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_728; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_729; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_730; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_731; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_732; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_733; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_734; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_735; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_736; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_737; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_738; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_739; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_740; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_741; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_742; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_743; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_744; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_745; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_746; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_747; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_748; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_749; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_750; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_751; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_752; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_753; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_754; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_755; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_756; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_757; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_758; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_759; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_760; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_761; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_762; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_763; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_764; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_765; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_766; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_767; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_768; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_769; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_770; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_771; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_772; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_773; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_774; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_775; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_776; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_777; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_778; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_779; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_780; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_781; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_782; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_783; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_784; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_785; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_786; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_787; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_788; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_789; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_790; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_791; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_792; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_793; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_794; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_795; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_796; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_797; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_798; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_799; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_800; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_801; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_802; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_803; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_804; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_805; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_806; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_807; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_808; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_809; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_810; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_811; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_812; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_813; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_814; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_815; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_816; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_817; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_818; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_819; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_820; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_821; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_822; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_823; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_824; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_825; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_826; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_827; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_828; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_829; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_830; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_831; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_832; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_833; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_834; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_835; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_836; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_837; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_838; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_839; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_840; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_841; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_842; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_843; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_844; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_845; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_846; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_847; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_848; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_849; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_850; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_851; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_852; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_853; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_854; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_855; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_856; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_857; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_858; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_859; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_860; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_861; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_862; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_863; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_864; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_865; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_866; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_867; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_868; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_869; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_870; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_871; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_872; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_873; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_874; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_875; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_876; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_877; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_878; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_879; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_880; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_881; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_882; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_883; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_884; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_885; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_886; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_887; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_888; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_889; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_890; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_891; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_892; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_893; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_894; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_895; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_896; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_897; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_898; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_899; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_900; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_901; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_902; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_903; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_904; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_905; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_906; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_907; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_908; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_909; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_910; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_911; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_912; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_913; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_914; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_915; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_916; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_917; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_918; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_919; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_920; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_921; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_922; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_923; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_924; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_925; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_926; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_927; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_928; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_929; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_930; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_931; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_932; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_933; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_934; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_935; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_936; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_937; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_938; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_939; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_940; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_941; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_942; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_943; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_944; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_945; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_946; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_947; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_948; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_949; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_950; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_951; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_952; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_953; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_954; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_955; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_956; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_957; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_958; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_959; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_960; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_961; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_962; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_963; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_964; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_965; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_966; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_967; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_968; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_969; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_970; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_971; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_972; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_973; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_974; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_975; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_976; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_977; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_978; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_979; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_980; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_981; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_982; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_983; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_984; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_985; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_986; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_987; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_988; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_989; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_990; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_991; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_992; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_993; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_994; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_995; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_996; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_997; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_998; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_999; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1000; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1001; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1002; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1003; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1004; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1005; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1006; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1007; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1008; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1009; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1010; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1011; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1012; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1013; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1014; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1015; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1016; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1017; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1018; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1019; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1020; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1021; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1022; // @[DataMemoryTest.scala 16:20]
  reg [31:0] mem_1023; // @[DataMemoryTest.scala 16:20]
  reg [31:0] io_dataOut_REG; // @[DataMemoryTest.scala 19:24]
  wire [31:0] _GEN_1 = 10'h1 == io_addr ? mem_1 : mem_0; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_2 = 10'h2 == io_addr ? mem_2 : _GEN_1; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_3 = 10'h3 == io_addr ? mem_3 : _GEN_2; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_4 = 10'h4 == io_addr ? mem_4 : _GEN_3; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_5 = 10'h5 == io_addr ? mem_5 : _GEN_4; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_6 = 10'h6 == io_addr ? mem_6 : _GEN_5; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_7 = 10'h7 == io_addr ? mem_7 : _GEN_6; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_8 = 10'h8 == io_addr ? mem_8 : _GEN_7; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_9 = 10'h9 == io_addr ? mem_9 : _GEN_8; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_10 = 10'ha == io_addr ? mem_10 : _GEN_9; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_11 = 10'hb == io_addr ? mem_11 : _GEN_10; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_12 = 10'hc == io_addr ? mem_12 : _GEN_11; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_13 = 10'hd == io_addr ? mem_13 : _GEN_12; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_14 = 10'he == io_addr ? mem_14 : _GEN_13; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_15 = 10'hf == io_addr ? mem_15 : _GEN_14; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_16 = 10'h10 == io_addr ? mem_16 : _GEN_15; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_17 = 10'h11 == io_addr ? mem_17 : _GEN_16; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_18 = 10'h12 == io_addr ? mem_18 : _GEN_17; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_19 = 10'h13 == io_addr ? mem_19 : _GEN_18; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_20 = 10'h14 == io_addr ? mem_20 : _GEN_19; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_21 = 10'h15 == io_addr ? mem_21 : _GEN_20; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_22 = 10'h16 == io_addr ? mem_22 : _GEN_21; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_23 = 10'h17 == io_addr ? mem_23 : _GEN_22; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_24 = 10'h18 == io_addr ? mem_24 : _GEN_23; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_25 = 10'h19 == io_addr ? mem_25 : _GEN_24; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_26 = 10'h1a == io_addr ? mem_26 : _GEN_25; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_27 = 10'h1b == io_addr ? mem_27 : _GEN_26; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_28 = 10'h1c == io_addr ? mem_28 : _GEN_27; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_29 = 10'h1d == io_addr ? mem_29 : _GEN_28; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_30 = 10'h1e == io_addr ? mem_30 : _GEN_29; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_31 = 10'h1f == io_addr ? mem_31 : _GEN_30; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_32 = 10'h20 == io_addr ? mem_32 : _GEN_31; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_33 = 10'h21 == io_addr ? mem_33 : _GEN_32; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_34 = 10'h22 == io_addr ? mem_34 : _GEN_33; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_35 = 10'h23 == io_addr ? mem_35 : _GEN_34; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_36 = 10'h24 == io_addr ? mem_36 : _GEN_35; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_37 = 10'h25 == io_addr ? mem_37 : _GEN_36; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_38 = 10'h26 == io_addr ? mem_38 : _GEN_37; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_39 = 10'h27 == io_addr ? mem_39 : _GEN_38; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_40 = 10'h28 == io_addr ? mem_40 : _GEN_39; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_41 = 10'h29 == io_addr ? mem_41 : _GEN_40; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_42 = 10'h2a == io_addr ? mem_42 : _GEN_41; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_43 = 10'h2b == io_addr ? mem_43 : _GEN_42; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_44 = 10'h2c == io_addr ? mem_44 : _GEN_43; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_45 = 10'h2d == io_addr ? mem_45 : _GEN_44; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_46 = 10'h2e == io_addr ? mem_46 : _GEN_45; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_47 = 10'h2f == io_addr ? mem_47 : _GEN_46; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_48 = 10'h30 == io_addr ? mem_48 : _GEN_47; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_49 = 10'h31 == io_addr ? mem_49 : _GEN_48; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_50 = 10'h32 == io_addr ? mem_50 : _GEN_49; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_51 = 10'h33 == io_addr ? mem_51 : _GEN_50; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_52 = 10'h34 == io_addr ? mem_52 : _GEN_51; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_53 = 10'h35 == io_addr ? mem_53 : _GEN_52; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_54 = 10'h36 == io_addr ? mem_54 : _GEN_53; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_55 = 10'h37 == io_addr ? mem_55 : _GEN_54; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_56 = 10'h38 == io_addr ? mem_56 : _GEN_55; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_57 = 10'h39 == io_addr ? mem_57 : _GEN_56; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_58 = 10'h3a == io_addr ? mem_58 : _GEN_57; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_59 = 10'h3b == io_addr ? mem_59 : _GEN_58; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_60 = 10'h3c == io_addr ? mem_60 : _GEN_59; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_61 = 10'h3d == io_addr ? mem_61 : _GEN_60; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_62 = 10'h3e == io_addr ? mem_62 : _GEN_61; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_63 = 10'h3f == io_addr ? mem_63 : _GEN_62; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_64 = 10'h40 == io_addr ? mem_64 : _GEN_63; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_65 = 10'h41 == io_addr ? mem_65 : _GEN_64; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_66 = 10'h42 == io_addr ? mem_66 : _GEN_65; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_67 = 10'h43 == io_addr ? mem_67 : _GEN_66; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_68 = 10'h44 == io_addr ? mem_68 : _GEN_67; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_69 = 10'h45 == io_addr ? mem_69 : _GEN_68; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_70 = 10'h46 == io_addr ? mem_70 : _GEN_69; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_71 = 10'h47 == io_addr ? mem_71 : _GEN_70; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_72 = 10'h48 == io_addr ? mem_72 : _GEN_71; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_73 = 10'h49 == io_addr ? mem_73 : _GEN_72; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_74 = 10'h4a == io_addr ? mem_74 : _GEN_73; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_75 = 10'h4b == io_addr ? mem_75 : _GEN_74; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_76 = 10'h4c == io_addr ? mem_76 : _GEN_75; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_77 = 10'h4d == io_addr ? mem_77 : _GEN_76; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_78 = 10'h4e == io_addr ? mem_78 : _GEN_77; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_79 = 10'h4f == io_addr ? mem_79 : _GEN_78; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_80 = 10'h50 == io_addr ? mem_80 : _GEN_79; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_81 = 10'h51 == io_addr ? mem_81 : _GEN_80; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_82 = 10'h52 == io_addr ? mem_82 : _GEN_81; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_83 = 10'h53 == io_addr ? mem_83 : _GEN_82; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_84 = 10'h54 == io_addr ? mem_84 : _GEN_83; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_85 = 10'h55 == io_addr ? mem_85 : _GEN_84; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_86 = 10'h56 == io_addr ? mem_86 : _GEN_85; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_87 = 10'h57 == io_addr ? mem_87 : _GEN_86; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_88 = 10'h58 == io_addr ? mem_88 : _GEN_87; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_89 = 10'h59 == io_addr ? mem_89 : _GEN_88; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_90 = 10'h5a == io_addr ? mem_90 : _GEN_89; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_91 = 10'h5b == io_addr ? mem_91 : _GEN_90; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_92 = 10'h5c == io_addr ? mem_92 : _GEN_91; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_93 = 10'h5d == io_addr ? mem_93 : _GEN_92; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_94 = 10'h5e == io_addr ? mem_94 : _GEN_93; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_95 = 10'h5f == io_addr ? mem_95 : _GEN_94; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_96 = 10'h60 == io_addr ? mem_96 : _GEN_95; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_97 = 10'h61 == io_addr ? mem_97 : _GEN_96; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_98 = 10'h62 == io_addr ? mem_98 : _GEN_97; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_99 = 10'h63 == io_addr ? mem_99 : _GEN_98; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_100 = 10'h64 == io_addr ? mem_100 : _GEN_99; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_101 = 10'h65 == io_addr ? mem_101 : _GEN_100; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_102 = 10'h66 == io_addr ? mem_102 : _GEN_101; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_103 = 10'h67 == io_addr ? mem_103 : _GEN_102; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_104 = 10'h68 == io_addr ? mem_104 : _GEN_103; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_105 = 10'h69 == io_addr ? mem_105 : _GEN_104; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_106 = 10'h6a == io_addr ? mem_106 : _GEN_105; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_107 = 10'h6b == io_addr ? mem_107 : _GEN_106; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_108 = 10'h6c == io_addr ? mem_108 : _GEN_107; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_109 = 10'h6d == io_addr ? mem_109 : _GEN_108; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_110 = 10'h6e == io_addr ? mem_110 : _GEN_109; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_111 = 10'h6f == io_addr ? mem_111 : _GEN_110; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_112 = 10'h70 == io_addr ? mem_112 : _GEN_111; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_113 = 10'h71 == io_addr ? mem_113 : _GEN_112; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_114 = 10'h72 == io_addr ? mem_114 : _GEN_113; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_115 = 10'h73 == io_addr ? mem_115 : _GEN_114; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_116 = 10'h74 == io_addr ? mem_116 : _GEN_115; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_117 = 10'h75 == io_addr ? mem_117 : _GEN_116; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_118 = 10'h76 == io_addr ? mem_118 : _GEN_117; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_119 = 10'h77 == io_addr ? mem_119 : _GEN_118; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_120 = 10'h78 == io_addr ? mem_120 : _GEN_119; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_121 = 10'h79 == io_addr ? mem_121 : _GEN_120; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_122 = 10'h7a == io_addr ? mem_122 : _GEN_121; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_123 = 10'h7b == io_addr ? mem_123 : _GEN_122; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_124 = 10'h7c == io_addr ? mem_124 : _GEN_123; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_125 = 10'h7d == io_addr ? mem_125 : _GEN_124; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_126 = 10'h7e == io_addr ? mem_126 : _GEN_125; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_127 = 10'h7f == io_addr ? mem_127 : _GEN_126; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_128 = 10'h80 == io_addr ? mem_128 : _GEN_127; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_129 = 10'h81 == io_addr ? mem_129 : _GEN_128; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_130 = 10'h82 == io_addr ? mem_130 : _GEN_129; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_131 = 10'h83 == io_addr ? mem_131 : _GEN_130; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_132 = 10'h84 == io_addr ? mem_132 : _GEN_131; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_133 = 10'h85 == io_addr ? mem_133 : _GEN_132; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_134 = 10'h86 == io_addr ? mem_134 : _GEN_133; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_135 = 10'h87 == io_addr ? mem_135 : _GEN_134; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_136 = 10'h88 == io_addr ? mem_136 : _GEN_135; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_137 = 10'h89 == io_addr ? mem_137 : _GEN_136; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_138 = 10'h8a == io_addr ? mem_138 : _GEN_137; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_139 = 10'h8b == io_addr ? mem_139 : _GEN_138; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_140 = 10'h8c == io_addr ? mem_140 : _GEN_139; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_141 = 10'h8d == io_addr ? mem_141 : _GEN_140; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_142 = 10'h8e == io_addr ? mem_142 : _GEN_141; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_143 = 10'h8f == io_addr ? mem_143 : _GEN_142; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_144 = 10'h90 == io_addr ? mem_144 : _GEN_143; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_145 = 10'h91 == io_addr ? mem_145 : _GEN_144; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_146 = 10'h92 == io_addr ? mem_146 : _GEN_145; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_147 = 10'h93 == io_addr ? mem_147 : _GEN_146; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_148 = 10'h94 == io_addr ? mem_148 : _GEN_147; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_149 = 10'h95 == io_addr ? mem_149 : _GEN_148; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_150 = 10'h96 == io_addr ? mem_150 : _GEN_149; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_151 = 10'h97 == io_addr ? mem_151 : _GEN_150; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_152 = 10'h98 == io_addr ? mem_152 : _GEN_151; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_153 = 10'h99 == io_addr ? mem_153 : _GEN_152; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_154 = 10'h9a == io_addr ? mem_154 : _GEN_153; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_155 = 10'h9b == io_addr ? mem_155 : _GEN_154; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_156 = 10'h9c == io_addr ? mem_156 : _GEN_155; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_157 = 10'h9d == io_addr ? mem_157 : _GEN_156; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_158 = 10'h9e == io_addr ? mem_158 : _GEN_157; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_159 = 10'h9f == io_addr ? mem_159 : _GEN_158; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_160 = 10'ha0 == io_addr ? mem_160 : _GEN_159; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_161 = 10'ha1 == io_addr ? mem_161 : _GEN_160; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_162 = 10'ha2 == io_addr ? mem_162 : _GEN_161; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_163 = 10'ha3 == io_addr ? mem_163 : _GEN_162; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_164 = 10'ha4 == io_addr ? mem_164 : _GEN_163; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_165 = 10'ha5 == io_addr ? mem_165 : _GEN_164; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_166 = 10'ha6 == io_addr ? mem_166 : _GEN_165; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_167 = 10'ha7 == io_addr ? mem_167 : _GEN_166; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_168 = 10'ha8 == io_addr ? mem_168 : _GEN_167; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_169 = 10'ha9 == io_addr ? mem_169 : _GEN_168; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_170 = 10'haa == io_addr ? mem_170 : _GEN_169; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_171 = 10'hab == io_addr ? mem_171 : _GEN_170; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_172 = 10'hac == io_addr ? mem_172 : _GEN_171; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_173 = 10'had == io_addr ? mem_173 : _GEN_172; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_174 = 10'hae == io_addr ? mem_174 : _GEN_173; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_175 = 10'haf == io_addr ? mem_175 : _GEN_174; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_176 = 10'hb0 == io_addr ? mem_176 : _GEN_175; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_177 = 10'hb1 == io_addr ? mem_177 : _GEN_176; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_178 = 10'hb2 == io_addr ? mem_178 : _GEN_177; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_179 = 10'hb3 == io_addr ? mem_179 : _GEN_178; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_180 = 10'hb4 == io_addr ? mem_180 : _GEN_179; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_181 = 10'hb5 == io_addr ? mem_181 : _GEN_180; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_182 = 10'hb6 == io_addr ? mem_182 : _GEN_181; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_183 = 10'hb7 == io_addr ? mem_183 : _GEN_182; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_184 = 10'hb8 == io_addr ? mem_184 : _GEN_183; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_185 = 10'hb9 == io_addr ? mem_185 : _GEN_184; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_186 = 10'hba == io_addr ? mem_186 : _GEN_185; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_187 = 10'hbb == io_addr ? mem_187 : _GEN_186; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_188 = 10'hbc == io_addr ? mem_188 : _GEN_187; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_189 = 10'hbd == io_addr ? mem_189 : _GEN_188; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_190 = 10'hbe == io_addr ? mem_190 : _GEN_189; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_191 = 10'hbf == io_addr ? mem_191 : _GEN_190; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_192 = 10'hc0 == io_addr ? mem_192 : _GEN_191; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_193 = 10'hc1 == io_addr ? mem_193 : _GEN_192; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_194 = 10'hc2 == io_addr ? mem_194 : _GEN_193; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_195 = 10'hc3 == io_addr ? mem_195 : _GEN_194; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_196 = 10'hc4 == io_addr ? mem_196 : _GEN_195; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_197 = 10'hc5 == io_addr ? mem_197 : _GEN_196; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_198 = 10'hc6 == io_addr ? mem_198 : _GEN_197; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_199 = 10'hc7 == io_addr ? mem_199 : _GEN_198; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_200 = 10'hc8 == io_addr ? mem_200 : _GEN_199; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_201 = 10'hc9 == io_addr ? mem_201 : _GEN_200; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_202 = 10'hca == io_addr ? mem_202 : _GEN_201; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_203 = 10'hcb == io_addr ? mem_203 : _GEN_202; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_204 = 10'hcc == io_addr ? mem_204 : _GEN_203; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_205 = 10'hcd == io_addr ? mem_205 : _GEN_204; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_206 = 10'hce == io_addr ? mem_206 : _GEN_205; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_207 = 10'hcf == io_addr ? mem_207 : _GEN_206; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_208 = 10'hd0 == io_addr ? mem_208 : _GEN_207; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_209 = 10'hd1 == io_addr ? mem_209 : _GEN_208; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_210 = 10'hd2 == io_addr ? mem_210 : _GEN_209; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_211 = 10'hd3 == io_addr ? mem_211 : _GEN_210; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_212 = 10'hd4 == io_addr ? mem_212 : _GEN_211; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_213 = 10'hd5 == io_addr ? mem_213 : _GEN_212; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_214 = 10'hd6 == io_addr ? mem_214 : _GEN_213; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_215 = 10'hd7 == io_addr ? mem_215 : _GEN_214; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_216 = 10'hd8 == io_addr ? mem_216 : _GEN_215; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_217 = 10'hd9 == io_addr ? mem_217 : _GEN_216; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_218 = 10'hda == io_addr ? mem_218 : _GEN_217; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_219 = 10'hdb == io_addr ? mem_219 : _GEN_218; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_220 = 10'hdc == io_addr ? mem_220 : _GEN_219; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_221 = 10'hdd == io_addr ? mem_221 : _GEN_220; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_222 = 10'hde == io_addr ? mem_222 : _GEN_221; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_223 = 10'hdf == io_addr ? mem_223 : _GEN_222; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_224 = 10'he0 == io_addr ? mem_224 : _GEN_223; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_225 = 10'he1 == io_addr ? mem_225 : _GEN_224; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_226 = 10'he2 == io_addr ? mem_226 : _GEN_225; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_227 = 10'he3 == io_addr ? mem_227 : _GEN_226; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_228 = 10'he4 == io_addr ? mem_228 : _GEN_227; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_229 = 10'he5 == io_addr ? mem_229 : _GEN_228; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_230 = 10'he6 == io_addr ? mem_230 : _GEN_229; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_231 = 10'he7 == io_addr ? mem_231 : _GEN_230; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_232 = 10'he8 == io_addr ? mem_232 : _GEN_231; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_233 = 10'he9 == io_addr ? mem_233 : _GEN_232; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_234 = 10'hea == io_addr ? mem_234 : _GEN_233; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_235 = 10'heb == io_addr ? mem_235 : _GEN_234; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_236 = 10'hec == io_addr ? mem_236 : _GEN_235; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_237 = 10'hed == io_addr ? mem_237 : _GEN_236; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_238 = 10'hee == io_addr ? mem_238 : _GEN_237; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_239 = 10'hef == io_addr ? mem_239 : _GEN_238; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_240 = 10'hf0 == io_addr ? mem_240 : _GEN_239; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_241 = 10'hf1 == io_addr ? mem_241 : _GEN_240; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_242 = 10'hf2 == io_addr ? mem_242 : _GEN_241; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_243 = 10'hf3 == io_addr ? mem_243 : _GEN_242; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_244 = 10'hf4 == io_addr ? mem_244 : _GEN_243; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_245 = 10'hf5 == io_addr ? mem_245 : _GEN_244; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_246 = 10'hf6 == io_addr ? mem_246 : _GEN_245; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_247 = 10'hf7 == io_addr ? mem_247 : _GEN_246; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_248 = 10'hf8 == io_addr ? mem_248 : _GEN_247; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_249 = 10'hf9 == io_addr ? mem_249 : _GEN_248; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_250 = 10'hfa == io_addr ? mem_250 : _GEN_249; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_251 = 10'hfb == io_addr ? mem_251 : _GEN_250; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_252 = 10'hfc == io_addr ? mem_252 : _GEN_251; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_253 = 10'hfd == io_addr ? mem_253 : _GEN_252; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_254 = 10'hfe == io_addr ? mem_254 : _GEN_253; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_255 = 10'hff == io_addr ? mem_255 : _GEN_254; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_256 = 10'h100 == io_addr ? mem_256 : _GEN_255; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_257 = 10'h101 == io_addr ? mem_257 : _GEN_256; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_258 = 10'h102 == io_addr ? mem_258 : _GEN_257; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_259 = 10'h103 == io_addr ? mem_259 : _GEN_258; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_260 = 10'h104 == io_addr ? mem_260 : _GEN_259; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_261 = 10'h105 == io_addr ? mem_261 : _GEN_260; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_262 = 10'h106 == io_addr ? mem_262 : _GEN_261; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_263 = 10'h107 == io_addr ? mem_263 : _GEN_262; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_264 = 10'h108 == io_addr ? mem_264 : _GEN_263; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_265 = 10'h109 == io_addr ? mem_265 : _GEN_264; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_266 = 10'h10a == io_addr ? mem_266 : _GEN_265; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_267 = 10'h10b == io_addr ? mem_267 : _GEN_266; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_268 = 10'h10c == io_addr ? mem_268 : _GEN_267; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_269 = 10'h10d == io_addr ? mem_269 : _GEN_268; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_270 = 10'h10e == io_addr ? mem_270 : _GEN_269; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_271 = 10'h10f == io_addr ? mem_271 : _GEN_270; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_272 = 10'h110 == io_addr ? mem_272 : _GEN_271; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_273 = 10'h111 == io_addr ? mem_273 : _GEN_272; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_274 = 10'h112 == io_addr ? mem_274 : _GEN_273; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_275 = 10'h113 == io_addr ? mem_275 : _GEN_274; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_276 = 10'h114 == io_addr ? mem_276 : _GEN_275; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_277 = 10'h115 == io_addr ? mem_277 : _GEN_276; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_278 = 10'h116 == io_addr ? mem_278 : _GEN_277; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_279 = 10'h117 == io_addr ? mem_279 : _GEN_278; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_280 = 10'h118 == io_addr ? mem_280 : _GEN_279; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_281 = 10'h119 == io_addr ? mem_281 : _GEN_280; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_282 = 10'h11a == io_addr ? mem_282 : _GEN_281; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_283 = 10'h11b == io_addr ? mem_283 : _GEN_282; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_284 = 10'h11c == io_addr ? mem_284 : _GEN_283; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_285 = 10'h11d == io_addr ? mem_285 : _GEN_284; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_286 = 10'h11e == io_addr ? mem_286 : _GEN_285; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_287 = 10'h11f == io_addr ? mem_287 : _GEN_286; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_288 = 10'h120 == io_addr ? mem_288 : _GEN_287; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_289 = 10'h121 == io_addr ? mem_289 : _GEN_288; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_290 = 10'h122 == io_addr ? mem_290 : _GEN_289; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_291 = 10'h123 == io_addr ? mem_291 : _GEN_290; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_292 = 10'h124 == io_addr ? mem_292 : _GEN_291; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_293 = 10'h125 == io_addr ? mem_293 : _GEN_292; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_294 = 10'h126 == io_addr ? mem_294 : _GEN_293; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_295 = 10'h127 == io_addr ? mem_295 : _GEN_294; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_296 = 10'h128 == io_addr ? mem_296 : _GEN_295; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_297 = 10'h129 == io_addr ? mem_297 : _GEN_296; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_298 = 10'h12a == io_addr ? mem_298 : _GEN_297; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_299 = 10'h12b == io_addr ? mem_299 : _GEN_298; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_300 = 10'h12c == io_addr ? mem_300 : _GEN_299; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_301 = 10'h12d == io_addr ? mem_301 : _GEN_300; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_302 = 10'h12e == io_addr ? mem_302 : _GEN_301; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_303 = 10'h12f == io_addr ? mem_303 : _GEN_302; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_304 = 10'h130 == io_addr ? mem_304 : _GEN_303; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_305 = 10'h131 == io_addr ? mem_305 : _GEN_304; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_306 = 10'h132 == io_addr ? mem_306 : _GEN_305; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_307 = 10'h133 == io_addr ? mem_307 : _GEN_306; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_308 = 10'h134 == io_addr ? mem_308 : _GEN_307; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_309 = 10'h135 == io_addr ? mem_309 : _GEN_308; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_310 = 10'h136 == io_addr ? mem_310 : _GEN_309; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_311 = 10'h137 == io_addr ? mem_311 : _GEN_310; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_312 = 10'h138 == io_addr ? mem_312 : _GEN_311; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_313 = 10'h139 == io_addr ? mem_313 : _GEN_312; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_314 = 10'h13a == io_addr ? mem_314 : _GEN_313; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_315 = 10'h13b == io_addr ? mem_315 : _GEN_314; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_316 = 10'h13c == io_addr ? mem_316 : _GEN_315; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_317 = 10'h13d == io_addr ? mem_317 : _GEN_316; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_318 = 10'h13e == io_addr ? mem_318 : _GEN_317; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_319 = 10'h13f == io_addr ? mem_319 : _GEN_318; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_320 = 10'h140 == io_addr ? mem_320 : _GEN_319; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_321 = 10'h141 == io_addr ? mem_321 : _GEN_320; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_322 = 10'h142 == io_addr ? mem_322 : _GEN_321; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_323 = 10'h143 == io_addr ? mem_323 : _GEN_322; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_324 = 10'h144 == io_addr ? mem_324 : _GEN_323; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_325 = 10'h145 == io_addr ? mem_325 : _GEN_324; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_326 = 10'h146 == io_addr ? mem_326 : _GEN_325; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_327 = 10'h147 == io_addr ? mem_327 : _GEN_326; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_328 = 10'h148 == io_addr ? mem_328 : _GEN_327; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_329 = 10'h149 == io_addr ? mem_329 : _GEN_328; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_330 = 10'h14a == io_addr ? mem_330 : _GEN_329; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_331 = 10'h14b == io_addr ? mem_331 : _GEN_330; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_332 = 10'h14c == io_addr ? mem_332 : _GEN_331; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_333 = 10'h14d == io_addr ? mem_333 : _GEN_332; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_334 = 10'h14e == io_addr ? mem_334 : _GEN_333; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_335 = 10'h14f == io_addr ? mem_335 : _GEN_334; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_336 = 10'h150 == io_addr ? mem_336 : _GEN_335; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_337 = 10'h151 == io_addr ? mem_337 : _GEN_336; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_338 = 10'h152 == io_addr ? mem_338 : _GEN_337; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_339 = 10'h153 == io_addr ? mem_339 : _GEN_338; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_340 = 10'h154 == io_addr ? mem_340 : _GEN_339; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_341 = 10'h155 == io_addr ? mem_341 : _GEN_340; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_342 = 10'h156 == io_addr ? mem_342 : _GEN_341; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_343 = 10'h157 == io_addr ? mem_343 : _GEN_342; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_344 = 10'h158 == io_addr ? mem_344 : _GEN_343; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_345 = 10'h159 == io_addr ? mem_345 : _GEN_344; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_346 = 10'h15a == io_addr ? mem_346 : _GEN_345; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_347 = 10'h15b == io_addr ? mem_347 : _GEN_346; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_348 = 10'h15c == io_addr ? mem_348 : _GEN_347; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_349 = 10'h15d == io_addr ? mem_349 : _GEN_348; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_350 = 10'h15e == io_addr ? mem_350 : _GEN_349; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_351 = 10'h15f == io_addr ? mem_351 : _GEN_350; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_352 = 10'h160 == io_addr ? mem_352 : _GEN_351; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_353 = 10'h161 == io_addr ? mem_353 : _GEN_352; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_354 = 10'h162 == io_addr ? mem_354 : _GEN_353; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_355 = 10'h163 == io_addr ? mem_355 : _GEN_354; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_356 = 10'h164 == io_addr ? mem_356 : _GEN_355; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_357 = 10'h165 == io_addr ? mem_357 : _GEN_356; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_358 = 10'h166 == io_addr ? mem_358 : _GEN_357; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_359 = 10'h167 == io_addr ? mem_359 : _GEN_358; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_360 = 10'h168 == io_addr ? mem_360 : _GEN_359; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_361 = 10'h169 == io_addr ? mem_361 : _GEN_360; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_362 = 10'h16a == io_addr ? mem_362 : _GEN_361; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_363 = 10'h16b == io_addr ? mem_363 : _GEN_362; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_364 = 10'h16c == io_addr ? mem_364 : _GEN_363; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_365 = 10'h16d == io_addr ? mem_365 : _GEN_364; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_366 = 10'h16e == io_addr ? mem_366 : _GEN_365; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_367 = 10'h16f == io_addr ? mem_367 : _GEN_366; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_368 = 10'h170 == io_addr ? mem_368 : _GEN_367; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_369 = 10'h171 == io_addr ? mem_369 : _GEN_368; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_370 = 10'h172 == io_addr ? mem_370 : _GEN_369; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_371 = 10'h173 == io_addr ? mem_371 : _GEN_370; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_372 = 10'h174 == io_addr ? mem_372 : _GEN_371; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_373 = 10'h175 == io_addr ? mem_373 : _GEN_372; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_374 = 10'h176 == io_addr ? mem_374 : _GEN_373; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_375 = 10'h177 == io_addr ? mem_375 : _GEN_374; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_376 = 10'h178 == io_addr ? mem_376 : _GEN_375; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_377 = 10'h179 == io_addr ? mem_377 : _GEN_376; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_378 = 10'h17a == io_addr ? mem_378 : _GEN_377; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_379 = 10'h17b == io_addr ? mem_379 : _GEN_378; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_380 = 10'h17c == io_addr ? mem_380 : _GEN_379; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_381 = 10'h17d == io_addr ? mem_381 : _GEN_380; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_382 = 10'h17e == io_addr ? mem_382 : _GEN_381; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_383 = 10'h17f == io_addr ? mem_383 : _GEN_382; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_384 = 10'h180 == io_addr ? mem_384 : _GEN_383; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_385 = 10'h181 == io_addr ? mem_385 : _GEN_384; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_386 = 10'h182 == io_addr ? mem_386 : _GEN_385; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_387 = 10'h183 == io_addr ? mem_387 : _GEN_386; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_388 = 10'h184 == io_addr ? mem_388 : _GEN_387; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_389 = 10'h185 == io_addr ? mem_389 : _GEN_388; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_390 = 10'h186 == io_addr ? mem_390 : _GEN_389; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_391 = 10'h187 == io_addr ? mem_391 : _GEN_390; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_392 = 10'h188 == io_addr ? mem_392 : _GEN_391; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_393 = 10'h189 == io_addr ? mem_393 : _GEN_392; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_394 = 10'h18a == io_addr ? mem_394 : _GEN_393; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_395 = 10'h18b == io_addr ? mem_395 : _GEN_394; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_396 = 10'h18c == io_addr ? mem_396 : _GEN_395; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_397 = 10'h18d == io_addr ? mem_397 : _GEN_396; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_398 = 10'h18e == io_addr ? mem_398 : _GEN_397; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_399 = 10'h18f == io_addr ? mem_399 : _GEN_398; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_400 = 10'h190 == io_addr ? mem_400 : _GEN_399; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_401 = 10'h191 == io_addr ? mem_401 : _GEN_400; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_402 = 10'h192 == io_addr ? mem_402 : _GEN_401; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_403 = 10'h193 == io_addr ? mem_403 : _GEN_402; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_404 = 10'h194 == io_addr ? mem_404 : _GEN_403; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_405 = 10'h195 == io_addr ? mem_405 : _GEN_404; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_406 = 10'h196 == io_addr ? mem_406 : _GEN_405; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_407 = 10'h197 == io_addr ? mem_407 : _GEN_406; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_408 = 10'h198 == io_addr ? mem_408 : _GEN_407; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_409 = 10'h199 == io_addr ? mem_409 : _GEN_408; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_410 = 10'h19a == io_addr ? mem_410 : _GEN_409; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_411 = 10'h19b == io_addr ? mem_411 : _GEN_410; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_412 = 10'h19c == io_addr ? mem_412 : _GEN_411; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_413 = 10'h19d == io_addr ? mem_413 : _GEN_412; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_414 = 10'h19e == io_addr ? mem_414 : _GEN_413; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_415 = 10'h19f == io_addr ? mem_415 : _GEN_414; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_416 = 10'h1a0 == io_addr ? mem_416 : _GEN_415; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_417 = 10'h1a1 == io_addr ? mem_417 : _GEN_416; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_418 = 10'h1a2 == io_addr ? mem_418 : _GEN_417; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_419 = 10'h1a3 == io_addr ? mem_419 : _GEN_418; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_420 = 10'h1a4 == io_addr ? mem_420 : _GEN_419; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_421 = 10'h1a5 == io_addr ? mem_421 : _GEN_420; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_422 = 10'h1a6 == io_addr ? mem_422 : _GEN_421; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_423 = 10'h1a7 == io_addr ? mem_423 : _GEN_422; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_424 = 10'h1a8 == io_addr ? mem_424 : _GEN_423; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_425 = 10'h1a9 == io_addr ? mem_425 : _GEN_424; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_426 = 10'h1aa == io_addr ? mem_426 : _GEN_425; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_427 = 10'h1ab == io_addr ? mem_427 : _GEN_426; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_428 = 10'h1ac == io_addr ? mem_428 : _GEN_427; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_429 = 10'h1ad == io_addr ? mem_429 : _GEN_428; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_430 = 10'h1ae == io_addr ? mem_430 : _GEN_429; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_431 = 10'h1af == io_addr ? mem_431 : _GEN_430; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_432 = 10'h1b0 == io_addr ? mem_432 : _GEN_431; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_433 = 10'h1b1 == io_addr ? mem_433 : _GEN_432; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_434 = 10'h1b2 == io_addr ? mem_434 : _GEN_433; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_435 = 10'h1b3 == io_addr ? mem_435 : _GEN_434; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_436 = 10'h1b4 == io_addr ? mem_436 : _GEN_435; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_437 = 10'h1b5 == io_addr ? mem_437 : _GEN_436; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_438 = 10'h1b6 == io_addr ? mem_438 : _GEN_437; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_439 = 10'h1b7 == io_addr ? mem_439 : _GEN_438; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_440 = 10'h1b8 == io_addr ? mem_440 : _GEN_439; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_441 = 10'h1b9 == io_addr ? mem_441 : _GEN_440; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_442 = 10'h1ba == io_addr ? mem_442 : _GEN_441; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_443 = 10'h1bb == io_addr ? mem_443 : _GEN_442; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_444 = 10'h1bc == io_addr ? mem_444 : _GEN_443; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_445 = 10'h1bd == io_addr ? mem_445 : _GEN_444; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_446 = 10'h1be == io_addr ? mem_446 : _GEN_445; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_447 = 10'h1bf == io_addr ? mem_447 : _GEN_446; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_448 = 10'h1c0 == io_addr ? mem_448 : _GEN_447; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_449 = 10'h1c1 == io_addr ? mem_449 : _GEN_448; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_450 = 10'h1c2 == io_addr ? mem_450 : _GEN_449; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_451 = 10'h1c3 == io_addr ? mem_451 : _GEN_450; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_452 = 10'h1c4 == io_addr ? mem_452 : _GEN_451; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_453 = 10'h1c5 == io_addr ? mem_453 : _GEN_452; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_454 = 10'h1c6 == io_addr ? mem_454 : _GEN_453; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_455 = 10'h1c7 == io_addr ? mem_455 : _GEN_454; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_456 = 10'h1c8 == io_addr ? mem_456 : _GEN_455; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_457 = 10'h1c9 == io_addr ? mem_457 : _GEN_456; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_458 = 10'h1ca == io_addr ? mem_458 : _GEN_457; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_459 = 10'h1cb == io_addr ? mem_459 : _GEN_458; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_460 = 10'h1cc == io_addr ? mem_460 : _GEN_459; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_461 = 10'h1cd == io_addr ? mem_461 : _GEN_460; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_462 = 10'h1ce == io_addr ? mem_462 : _GEN_461; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_463 = 10'h1cf == io_addr ? mem_463 : _GEN_462; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_464 = 10'h1d0 == io_addr ? mem_464 : _GEN_463; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_465 = 10'h1d1 == io_addr ? mem_465 : _GEN_464; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_466 = 10'h1d2 == io_addr ? mem_466 : _GEN_465; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_467 = 10'h1d3 == io_addr ? mem_467 : _GEN_466; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_468 = 10'h1d4 == io_addr ? mem_468 : _GEN_467; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_469 = 10'h1d5 == io_addr ? mem_469 : _GEN_468; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_470 = 10'h1d6 == io_addr ? mem_470 : _GEN_469; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_471 = 10'h1d7 == io_addr ? mem_471 : _GEN_470; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_472 = 10'h1d8 == io_addr ? mem_472 : _GEN_471; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_473 = 10'h1d9 == io_addr ? mem_473 : _GEN_472; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_474 = 10'h1da == io_addr ? mem_474 : _GEN_473; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_475 = 10'h1db == io_addr ? mem_475 : _GEN_474; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_476 = 10'h1dc == io_addr ? mem_476 : _GEN_475; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_477 = 10'h1dd == io_addr ? mem_477 : _GEN_476; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_478 = 10'h1de == io_addr ? mem_478 : _GEN_477; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_479 = 10'h1df == io_addr ? mem_479 : _GEN_478; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_480 = 10'h1e0 == io_addr ? mem_480 : _GEN_479; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_481 = 10'h1e1 == io_addr ? mem_481 : _GEN_480; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_482 = 10'h1e2 == io_addr ? mem_482 : _GEN_481; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_483 = 10'h1e3 == io_addr ? mem_483 : _GEN_482; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_484 = 10'h1e4 == io_addr ? mem_484 : _GEN_483; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_485 = 10'h1e5 == io_addr ? mem_485 : _GEN_484; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_486 = 10'h1e6 == io_addr ? mem_486 : _GEN_485; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_487 = 10'h1e7 == io_addr ? mem_487 : _GEN_486; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_488 = 10'h1e8 == io_addr ? mem_488 : _GEN_487; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_489 = 10'h1e9 == io_addr ? mem_489 : _GEN_488; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_490 = 10'h1ea == io_addr ? mem_490 : _GEN_489; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_491 = 10'h1eb == io_addr ? mem_491 : _GEN_490; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_492 = 10'h1ec == io_addr ? mem_492 : _GEN_491; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_493 = 10'h1ed == io_addr ? mem_493 : _GEN_492; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_494 = 10'h1ee == io_addr ? mem_494 : _GEN_493; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_495 = 10'h1ef == io_addr ? mem_495 : _GEN_494; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_496 = 10'h1f0 == io_addr ? mem_496 : _GEN_495; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_497 = 10'h1f1 == io_addr ? mem_497 : _GEN_496; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_498 = 10'h1f2 == io_addr ? mem_498 : _GEN_497; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_499 = 10'h1f3 == io_addr ? mem_499 : _GEN_498; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_500 = 10'h1f4 == io_addr ? mem_500 : _GEN_499; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_501 = 10'h1f5 == io_addr ? mem_501 : _GEN_500; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_502 = 10'h1f6 == io_addr ? mem_502 : _GEN_501; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_503 = 10'h1f7 == io_addr ? mem_503 : _GEN_502; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_504 = 10'h1f8 == io_addr ? mem_504 : _GEN_503; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_505 = 10'h1f9 == io_addr ? mem_505 : _GEN_504; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_506 = 10'h1fa == io_addr ? mem_506 : _GEN_505; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_507 = 10'h1fb == io_addr ? mem_507 : _GEN_506; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_508 = 10'h1fc == io_addr ? mem_508 : _GEN_507; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_509 = 10'h1fd == io_addr ? mem_509 : _GEN_508; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_510 = 10'h1fe == io_addr ? mem_510 : _GEN_509; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_511 = 10'h1ff == io_addr ? mem_511 : _GEN_510; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_512 = 10'h200 == io_addr ? mem_512 : _GEN_511; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_513 = 10'h201 == io_addr ? mem_513 : _GEN_512; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_514 = 10'h202 == io_addr ? mem_514 : _GEN_513; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_515 = 10'h203 == io_addr ? mem_515 : _GEN_514; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_516 = 10'h204 == io_addr ? mem_516 : _GEN_515; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_517 = 10'h205 == io_addr ? mem_517 : _GEN_516; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_518 = 10'h206 == io_addr ? mem_518 : _GEN_517; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_519 = 10'h207 == io_addr ? mem_519 : _GEN_518; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_520 = 10'h208 == io_addr ? mem_520 : _GEN_519; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_521 = 10'h209 == io_addr ? mem_521 : _GEN_520; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_522 = 10'h20a == io_addr ? mem_522 : _GEN_521; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_523 = 10'h20b == io_addr ? mem_523 : _GEN_522; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_524 = 10'h20c == io_addr ? mem_524 : _GEN_523; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_525 = 10'h20d == io_addr ? mem_525 : _GEN_524; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_526 = 10'h20e == io_addr ? mem_526 : _GEN_525; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_527 = 10'h20f == io_addr ? mem_527 : _GEN_526; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_528 = 10'h210 == io_addr ? mem_528 : _GEN_527; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_529 = 10'h211 == io_addr ? mem_529 : _GEN_528; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_530 = 10'h212 == io_addr ? mem_530 : _GEN_529; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_531 = 10'h213 == io_addr ? mem_531 : _GEN_530; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_532 = 10'h214 == io_addr ? mem_532 : _GEN_531; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_533 = 10'h215 == io_addr ? mem_533 : _GEN_532; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_534 = 10'h216 == io_addr ? mem_534 : _GEN_533; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_535 = 10'h217 == io_addr ? mem_535 : _GEN_534; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_536 = 10'h218 == io_addr ? mem_536 : _GEN_535; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_537 = 10'h219 == io_addr ? mem_537 : _GEN_536; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_538 = 10'h21a == io_addr ? mem_538 : _GEN_537; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_539 = 10'h21b == io_addr ? mem_539 : _GEN_538; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_540 = 10'h21c == io_addr ? mem_540 : _GEN_539; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_541 = 10'h21d == io_addr ? mem_541 : _GEN_540; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_542 = 10'h21e == io_addr ? mem_542 : _GEN_541; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_543 = 10'h21f == io_addr ? mem_543 : _GEN_542; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_544 = 10'h220 == io_addr ? mem_544 : _GEN_543; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_545 = 10'h221 == io_addr ? mem_545 : _GEN_544; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_546 = 10'h222 == io_addr ? mem_546 : _GEN_545; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_547 = 10'h223 == io_addr ? mem_547 : _GEN_546; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_548 = 10'h224 == io_addr ? mem_548 : _GEN_547; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_549 = 10'h225 == io_addr ? mem_549 : _GEN_548; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_550 = 10'h226 == io_addr ? mem_550 : _GEN_549; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_551 = 10'h227 == io_addr ? mem_551 : _GEN_550; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_552 = 10'h228 == io_addr ? mem_552 : _GEN_551; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_553 = 10'h229 == io_addr ? mem_553 : _GEN_552; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_554 = 10'h22a == io_addr ? mem_554 : _GEN_553; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_555 = 10'h22b == io_addr ? mem_555 : _GEN_554; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_556 = 10'h22c == io_addr ? mem_556 : _GEN_555; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_557 = 10'h22d == io_addr ? mem_557 : _GEN_556; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_558 = 10'h22e == io_addr ? mem_558 : _GEN_557; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_559 = 10'h22f == io_addr ? mem_559 : _GEN_558; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_560 = 10'h230 == io_addr ? mem_560 : _GEN_559; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_561 = 10'h231 == io_addr ? mem_561 : _GEN_560; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_562 = 10'h232 == io_addr ? mem_562 : _GEN_561; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_563 = 10'h233 == io_addr ? mem_563 : _GEN_562; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_564 = 10'h234 == io_addr ? mem_564 : _GEN_563; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_565 = 10'h235 == io_addr ? mem_565 : _GEN_564; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_566 = 10'h236 == io_addr ? mem_566 : _GEN_565; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_567 = 10'h237 == io_addr ? mem_567 : _GEN_566; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_568 = 10'h238 == io_addr ? mem_568 : _GEN_567; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_569 = 10'h239 == io_addr ? mem_569 : _GEN_568; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_570 = 10'h23a == io_addr ? mem_570 : _GEN_569; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_571 = 10'h23b == io_addr ? mem_571 : _GEN_570; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_572 = 10'h23c == io_addr ? mem_572 : _GEN_571; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_573 = 10'h23d == io_addr ? mem_573 : _GEN_572; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_574 = 10'h23e == io_addr ? mem_574 : _GEN_573; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_575 = 10'h23f == io_addr ? mem_575 : _GEN_574; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_576 = 10'h240 == io_addr ? mem_576 : _GEN_575; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_577 = 10'h241 == io_addr ? mem_577 : _GEN_576; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_578 = 10'h242 == io_addr ? mem_578 : _GEN_577; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_579 = 10'h243 == io_addr ? mem_579 : _GEN_578; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_580 = 10'h244 == io_addr ? mem_580 : _GEN_579; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_581 = 10'h245 == io_addr ? mem_581 : _GEN_580; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_582 = 10'h246 == io_addr ? mem_582 : _GEN_581; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_583 = 10'h247 == io_addr ? mem_583 : _GEN_582; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_584 = 10'h248 == io_addr ? mem_584 : _GEN_583; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_585 = 10'h249 == io_addr ? mem_585 : _GEN_584; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_586 = 10'h24a == io_addr ? mem_586 : _GEN_585; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_587 = 10'h24b == io_addr ? mem_587 : _GEN_586; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_588 = 10'h24c == io_addr ? mem_588 : _GEN_587; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_589 = 10'h24d == io_addr ? mem_589 : _GEN_588; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_590 = 10'h24e == io_addr ? mem_590 : _GEN_589; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_591 = 10'h24f == io_addr ? mem_591 : _GEN_590; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_592 = 10'h250 == io_addr ? mem_592 : _GEN_591; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_593 = 10'h251 == io_addr ? mem_593 : _GEN_592; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_594 = 10'h252 == io_addr ? mem_594 : _GEN_593; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_595 = 10'h253 == io_addr ? mem_595 : _GEN_594; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_596 = 10'h254 == io_addr ? mem_596 : _GEN_595; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_597 = 10'h255 == io_addr ? mem_597 : _GEN_596; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_598 = 10'h256 == io_addr ? mem_598 : _GEN_597; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_599 = 10'h257 == io_addr ? mem_599 : _GEN_598; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_600 = 10'h258 == io_addr ? mem_600 : _GEN_599; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_601 = 10'h259 == io_addr ? mem_601 : _GEN_600; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_602 = 10'h25a == io_addr ? mem_602 : _GEN_601; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_603 = 10'h25b == io_addr ? mem_603 : _GEN_602; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_604 = 10'h25c == io_addr ? mem_604 : _GEN_603; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_605 = 10'h25d == io_addr ? mem_605 : _GEN_604; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_606 = 10'h25e == io_addr ? mem_606 : _GEN_605; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_607 = 10'h25f == io_addr ? mem_607 : _GEN_606; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_608 = 10'h260 == io_addr ? mem_608 : _GEN_607; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_609 = 10'h261 == io_addr ? mem_609 : _GEN_608; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_610 = 10'h262 == io_addr ? mem_610 : _GEN_609; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_611 = 10'h263 == io_addr ? mem_611 : _GEN_610; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_612 = 10'h264 == io_addr ? mem_612 : _GEN_611; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_613 = 10'h265 == io_addr ? mem_613 : _GEN_612; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_614 = 10'h266 == io_addr ? mem_614 : _GEN_613; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_615 = 10'h267 == io_addr ? mem_615 : _GEN_614; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_616 = 10'h268 == io_addr ? mem_616 : _GEN_615; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_617 = 10'h269 == io_addr ? mem_617 : _GEN_616; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_618 = 10'h26a == io_addr ? mem_618 : _GEN_617; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_619 = 10'h26b == io_addr ? mem_619 : _GEN_618; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_620 = 10'h26c == io_addr ? mem_620 : _GEN_619; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_621 = 10'h26d == io_addr ? mem_621 : _GEN_620; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_622 = 10'h26e == io_addr ? mem_622 : _GEN_621; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_623 = 10'h26f == io_addr ? mem_623 : _GEN_622; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_624 = 10'h270 == io_addr ? mem_624 : _GEN_623; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_625 = 10'h271 == io_addr ? mem_625 : _GEN_624; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_626 = 10'h272 == io_addr ? mem_626 : _GEN_625; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_627 = 10'h273 == io_addr ? mem_627 : _GEN_626; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_628 = 10'h274 == io_addr ? mem_628 : _GEN_627; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_629 = 10'h275 == io_addr ? mem_629 : _GEN_628; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_630 = 10'h276 == io_addr ? mem_630 : _GEN_629; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_631 = 10'h277 == io_addr ? mem_631 : _GEN_630; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_632 = 10'h278 == io_addr ? mem_632 : _GEN_631; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_633 = 10'h279 == io_addr ? mem_633 : _GEN_632; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_634 = 10'h27a == io_addr ? mem_634 : _GEN_633; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_635 = 10'h27b == io_addr ? mem_635 : _GEN_634; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_636 = 10'h27c == io_addr ? mem_636 : _GEN_635; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_637 = 10'h27d == io_addr ? mem_637 : _GEN_636; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_638 = 10'h27e == io_addr ? mem_638 : _GEN_637; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_639 = 10'h27f == io_addr ? mem_639 : _GEN_638; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_640 = 10'h280 == io_addr ? mem_640 : _GEN_639; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_641 = 10'h281 == io_addr ? mem_641 : _GEN_640; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_642 = 10'h282 == io_addr ? mem_642 : _GEN_641; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_643 = 10'h283 == io_addr ? mem_643 : _GEN_642; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_644 = 10'h284 == io_addr ? mem_644 : _GEN_643; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_645 = 10'h285 == io_addr ? mem_645 : _GEN_644; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_646 = 10'h286 == io_addr ? mem_646 : _GEN_645; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_647 = 10'h287 == io_addr ? mem_647 : _GEN_646; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_648 = 10'h288 == io_addr ? mem_648 : _GEN_647; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_649 = 10'h289 == io_addr ? mem_649 : _GEN_648; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_650 = 10'h28a == io_addr ? mem_650 : _GEN_649; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_651 = 10'h28b == io_addr ? mem_651 : _GEN_650; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_652 = 10'h28c == io_addr ? mem_652 : _GEN_651; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_653 = 10'h28d == io_addr ? mem_653 : _GEN_652; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_654 = 10'h28e == io_addr ? mem_654 : _GEN_653; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_655 = 10'h28f == io_addr ? mem_655 : _GEN_654; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_656 = 10'h290 == io_addr ? mem_656 : _GEN_655; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_657 = 10'h291 == io_addr ? mem_657 : _GEN_656; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_658 = 10'h292 == io_addr ? mem_658 : _GEN_657; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_659 = 10'h293 == io_addr ? mem_659 : _GEN_658; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_660 = 10'h294 == io_addr ? mem_660 : _GEN_659; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_661 = 10'h295 == io_addr ? mem_661 : _GEN_660; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_662 = 10'h296 == io_addr ? mem_662 : _GEN_661; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_663 = 10'h297 == io_addr ? mem_663 : _GEN_662; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_664 = 10'h298 == io_addr ? mem_664 : _GEN_663; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_665 = 10'h299 == io_addr ? mem_665 : _GEN_664; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_666 = 10'h29a == io_addr ? mem_666 : _GEN_665; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_667 = 10'h29b == io_addr ? mem_667 : _GEN_666; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_668 = 10'h29c == io_addr ? mem_668 : _GEN_667; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_669 = 10'h29d == io_addr ? mem_669 : _GEN_668; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_670 = 10'h29e == io_addr ? mem_670 : _GEN_669; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_671 = 10'h29f == io_addr ? mem_671 : _GEN_670; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_672 = 10'h2a0 == io_addr ? mem_672 : _GEN_671; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_673 = 10'h2a1 == io_addr ? mem_673 : _GEN_672; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_674 = 10'h2a2 == io_addr ? mem_674 : _GEN_673; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_675 = 10'h2a3 == io_addr ? mem_675 : _GEN_674; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_676 = 10'h2a4 == io_addr ? mem_676 : _GEN_675; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_677 = 10'h2a5 == io_addr ? mem_677 : _GEN_676; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_678 = 10'h2a6 == io_addr ? mem_678 : _GEN_677; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_679 = 10'h2a7 == io_addr ? mem_679 : _GEN_678; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_680 = 10'h2a8 == io_addr ? mem_680 : _GEN_679; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_681 = 10'h2a9 == io_addr ? mem_681 : _GEN_680; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_682 = 10'h2aa == io_addr ? mem_682 : _GEN_681; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_683 = 10'h2ab == io_addr ? mem_683 : _GEN_682; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_684 = 10'h2ac == io_addr ? mem_684 : _GEN_683; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_685 = 10'h2ad == io_addr ? mem_685 : _GEN_684; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_686 = 10'h2ae == io_addr ? mem_686 : _GEN_685; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_687 = 10'h2af == io_addr ? mem_687 : _GEN_686; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_688 = 10'h2b0 == io_addr ? mem_688 : _GEN_687; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_689 = 10'h2b1 == io_addr ? mem_689 : _GEN_688; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_690 = 10'h2b2 == io_addr ? mem_690 : _GEN_689; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_691 = 10'h2b3 == io_addr ? mem_691 : _GEN_690; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_692 = 10'h2b4 == io_addr ? mem_692 : _GEN_691; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_693 = 10'h2b5 == io_addr ? mem_693 : _GEN_692; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_694 = 10'h2b6 == io_addr ? mem_694 : _GEN_693; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_695 = 10'h2b7 == io_addr ? mem_695 : _GEN_694; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_696 = 10'h2b8 == io_addr ? mem_696 : _GEN_695; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_697 = 10'h2b9 == io_addr ? mem_697 : _GEN_696; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_698 = 10'h2ba == io_addr ? mem_698 : _GEN_697; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_699 = 10'h2bb == io_addr ? mem_699 : _GEN_698; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_700 = 10'h2bc == io_addr ? mem_700 : _GEN_699; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_701 = 10'h2bd == io_addr ? mem_701 : _GEN_700; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_702 = 10'h2be == io_addr ? mem_702 : _GEN_701; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_703 = 10'h2bf == io_addr ? mem_703 : _GEN_702; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_704 = 10'h2c0 == io_addr ? mem_704 : _GEN_703; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_705 = 10'h2c1 == io_addr ? mem_705 : _GEN_704; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_706 = 10'h2c2 == io_addr ? mem_706 : _GEN_705; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_707 = 10'h2c3 == io_addr ? mem_707 : _GEN_706; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_708 = 10'h2c4 == io_addr ? mem_708 : _GEN_707; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_709 = 10'h2c5 == io_addr ? mem_709 : _GEN_708; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_710 = 10'h2c6 == io_addr ? mem_710 : _GEN_709; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_711 = 10'h2c7 == io_addr ? mem_711 : _GEN_710; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_712 = 10'h2c8 == io_addr ? mem_712 : _GEN_711; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_713 = 10'h2c9 == io_addr ? mem_713 : _GEN_712; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_714 = 10'h2ca == io_addr ? mem_714 : _GEN_713; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_715 = 10'h2cb == io_addr ? mem_715 : _GEN_714; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_716 = 10'h2cc == io_addr ? mem_716 : _GEN_715; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_717 = 10'h2cd == io_addr ? mem_717 : _GEN_716; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_718 = 10'h2ce == io_addr ? mem_718 : _GEN_717; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_719 = 10'h2cf == io_addr ? mem_719 : _GEN_718; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_720 = 10'h2d0 == io_addr ? mem_720 : _GEN_719; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_721 = 10'h2d1 == io_addr ? mem_721 : _GEN_720; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_722 = 10'h2d2 == io_addr ? mem_722 : _GEN_721; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_723 = 10'h2d3 == io_addr ? mem_723 : _GEN_722; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_724 = 10'h2d4 == io_addr ? mem_724 : _GEN_723; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_725 = 10'h2d5 == io_addr ? mem_725 : _GEN_724; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_726 = 10'h2d6 == io_addr ? mem_726 : _GEN_725; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_727 = 10'h2d7 == io_addr ? mem_727 : _GEN_726; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_728 = 10'h2d8 == io_addr ? mem_728 : _GEN_727; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_729 = 10'h2d9 == io_addr ? mem_729 : _GEN_728; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_730 = 10'h2da == io_addr ? mem_730 : _GEN_729; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_731 = 10'h2db == io_addr ? mem_731 : _GEN_730; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_732 = 10'h2dc == io_addr ? mem_732 : _GEN_731; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_733 = 10'h2dd == io_addr ? mem_733 : _GEN_732; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_734 = 10'h2de == io_addr ? mem_734 : _GEN_733; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_735 = 10'h2df == io_addr ? mem_735 : _GEN_734; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_736 = 10'h2e0 == io_addr ? mem_736 : _GEN_735; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_737 = 10'h2e1 == io_addr ? mem_737 : _GEN_736; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_738 = 10'h2e2 == io_addr ? mem_738 : _GEN_737; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_739 = 10'h2e3 == io_addr ? mem_739 : _GEN_738; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_740 = 10'h2e4 == io_addr ? mem_740 : _GEN_739; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_741 = 10'h2e5 == io_addr ? mem_741 : _GEN_740; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_742 = 10'h2e6 == io_addr ? mem_742 : _GEN_741; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_743 = 10'h2e7 == io_addr ? mem_743 : _GEN_742; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_744 = 10'h2e8 == io_addr ? mem_744 : _GEN_743; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_745 = 10'h2e9 == io_addr ? mem_745 : _GEN_744; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_746 = 10'h2ea == io_addr ? mem_746 : _GEN_745; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_747 = 10'h2eb == io_addr ? mem_747 : _GEN_746; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_748 = 10'h2ec == io_addr ? mem_748 : _GEN_747; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_749 = 10'h2ed == io_addr ? mem_749 : _GEN_748; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_750 = 10'h2ee == io_addr ? mem_750 : _GEN_749; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_751 = 10'h2ef == io_addr ? mem_751 : _GEN_750; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_752 = 10'h2f0 == io_addr ? mem_752 : _GEN_751; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_753 = 10'h2f1 == io_addr ? mem_753 : _GEN_752; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_754 = 10'h2f2 == io_addr ? mem_754 : _GEN_753; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_755 = 10'h2f3 == io_addr ? mem_755 : _GEN_754; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_756 = 10'h2f4 == io_addr ? mem_756 : _GEN_755; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_757 = 10'h2f5 == io_addr ? mem_757 : _GEN_756; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_758 = 10'h2f6 == io_addr ? mem_758 : _GEN_757; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_759 = 10'h2f7 == io_addr ? mem_759 : _GEN_758; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_760 = 10'h2f8 == io_addr ? mem_760 : _GEN_759; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_761 = 10'h2f9 == io_addr ? mem_761 : _GEN_760; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_762 = 10'h2fa == io_addr ? mem_762 : _GEN_761; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_763 = 10'h2fb == io_addr ? mem_763 : _GEN_762; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_764 = 10'h2fc == io_addr ? mem_764 : _GEN_763; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_765 = 10'h2fd == io_addr ? mem_765 : _GEN_764; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_766 = 10'h2fe == io_addr ? mem_766 : _GEN_765; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_767 = 10'h2ff == io_addr ? mem_767 : _GEN_766; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_768 = 10'h300 == io_addr ? mem_768 : _GEN_767; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_769 = 10'h301 == io_addr ? mem_769 : _GEN_768; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_770 = 10'h302 == io_addr ? mem_770 : _GEN_769; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_771 = 10'h303 == io_addr ? mem_771 : _GEN_770; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_772 = 10'h304 == io_addr ? mem_772 : _GEN_771; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_773 = 10'h305 == io_addr ? mem_773 : _GEN_772; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_774 = 10'h306 == io_addr ? mem_774 : _GEN_773; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_775 = 10'h307 == io_addr ? mem_775 : _GEN_774; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_776 = 10'h308 == io_addr ? mem_776 : _GEN_775; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_777 = 10'h309 == io_addr ? mem_777 : _GEN_776; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_778 = 10'h30a == io_addr ? mem_778 : _GEN_777; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_779 = 10'h30b == io_addr ? mem_779 : _GEN_778; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_780 = 10'h30c == io_addr ? mem_780 : _GEN_779; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_781 = 10'h30d == io_addr ? mem_781 : _GEN_780; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_782 = 10'h30e == io_addr ? mem_782 : _GEN_781; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_783 = 10'h30f == io_addr ? mem_783 : _GEN_782; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_784 = 10'h310 == io_addr ? mem_784 : _GEN_783; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_785 = 10'h311 == io_addr ? mem_785 : _GEN_784; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_786 = 10'h312 == io_addr ? mem_786 : _GEN_785; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_787 = 10'h313 == io_addr ? mem_787 : _GEN_786; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_788 = 10'h314 == io_addr ? mem_788 : _GEN_787; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_789 = 10'h315 == io_addr ? mem_789 : _GEN_788; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_790 = 10'h316 == io_addr ? mem_790 : _GEN_789; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_791 = 10'h317 == io_addr ? mem_791 : _GEN_790; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_792 = 10'h318 == io_addr ? mem_792 : _GEN_791; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_793 = 10'h319 == io_addr ? mem_793 : _GEN_792; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_794 = 10'h31a == io_addr ? mem_794 : _GEN_793; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_795 = 10'h31b == io_addr ? mem_795 : _GEN_794; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_796 = 10'h31c == io_addr ? mem_796 : _GEN_795; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_797 = 10'h31d == io_addr ? mem_797 : _GEN_796; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_798 = 10'h31e == io_addr ? mem_798 : _GEN_797; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_799 = 10'h31f == io_addr ? mem_799 : _GEN_798; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_800 = 10'h320 == io_addr ? mem_800 : _GEN_799; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_801 = 10'h321 == io_addr ? mem_801 : _GEN_800; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_802 = 10'h322 == io_addr ? mem_802 : _GEN_801; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_803 = 10'h323 == io_addr ? mem_803 : _GEN_802; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_804 = 10'h324 == io_addr ? mem_804 : _GEN_803; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_805 = 10'h325 == io_addr ? mem_805 : _GEN_804; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_806 = 10'h326 == io_addr ? mem_806 : _GEN_805; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_807 = 10'h327 == io_addr ? mem_807 : _GEN_806; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_808 = 10'h328 == io_addr ? mem_808 : _GEN_807; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_809 = 10'h329 == io_addr ? mem_809 : _GEN_808; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_810 = 10'h32a == io_addr ? mem_810 : _GEN_809; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_811 = 10'h32b == io_addr ? mem_811 : _GEN_810; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_812 = 10'h32c == io_addr ? mem_812 : _GEN_811; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_813 = 10'h32d == io_addr ? mem_813 : _GEN_812; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_814 = 10'h32e == io_addr ? mem_814 : _GEN_813; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_815 = 10'h32f == io_addr ? mem_815 : _GEN_814; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_816 = 10'h330 == io_addr ? mem_816 : _GEN_815; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_817 = 10'h331 == io_addr ? mem_817 : _GEN_816; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_818 = 10'h332 == io_addr ? mem_818 : _GEN_817; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_819 = 10'h333 == io_addr ? mem_819 : _GEN_818; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_820 = 10'h334 == io_addr ? mem_820 : _GEN_819; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_821 = 10'h335 == io_addr ? mem_821 : _GEN_820; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_822 = 10'h336 == io_addr ? mem_822 : _GEN_821; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_823 = 10'h337 == io_addr ? mem_823 : _GEN_822; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_824 = 10'h338 == io_addr ? mem_824 : _GEN_823; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_825 = 10'h339 == io_addr ? mem_825 : _GEN_824; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_826 = 10'h33a == io_addr ? mem_826 : _GEN_825; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_827 = 10'h33b == io_addr ? mem_827 : _GEN_826; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_828 = 10'h33c == io_addr ? mem_828 : _GEN_827; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_829 = 10'h33d == io_addr ? mem_829 : _GEN_828; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_830 = 10'h33e == io_addr ? mem_830 : _GEN_829; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_831 = 10'h33f == io_addr ? mem_831 : _GEN_830; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_832 = 10'h340 == io_addr ? mem_832 : _GEN_831; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_833 = 10'h341 == io_addr ? mem_833 : _GEN_832; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_834 = 10'h342 == io_addr ? mem_834 : _GEN_833; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_835 = 10'h343 == io_addr ? mem_835 : _GEN_834; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_836 = 10'h344 == io_addr ? mem_836 : _GEN_835; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_837 = 10'h345 == io_addr ? mem_837 : _GEN_836; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_838 = 10'h346 == io_addr ? mem_838 : _GEN_837; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_839 = 10'h347 == io_addr ? mem_839 : _GEN_838; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_840 = 10'h348 == io_addr ? mem_840 : _GEN_839; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_841 = 10'h349 == io_addr ? mem_841 : _GEN_840; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_842 = 10'h34a == io_addr ? mem_842 : _GEN_841; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_843 = 10'h34b == io_addr ? mem_843 : _GEN_842; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_844 = 10'h34c == io_addr ? mem_844 : _GEN_843; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_845 = 10'h34d == io_addr ? mem_845 : _GEN_844; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_846 = 10'h34e == io_addr ? mem_846 : _GEN_845; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_847 = 10'h34f == io_addr ? mem_847 : _GEN_846; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_848 = 10'h350 == io_addr ? mem_848 : _GEN_847; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_849 = 10'h351 == io_addr ? mem_849 : _GEN_848; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_850 = 10'h352 == io_addr ? mem_850 : _GEN_849; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_851 = 10'h353 == io_addr ? mem_851 : _GEN_850; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_852 = 10'h354 == io_addr ? mem_852 : _GEN_851; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_853 = 10'h355 == io_addr ? mem_853 : _GEN_852; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_854 = 10'h356 == io_addr ? mem_854 : _GEN_853; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_855 = 10'h357 == io_addr ? mem_855 : _GEN_854; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_856 = 10'h358 == io_addr ? mem_856 : _GEN_855; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_857 = 10'h359 == io_addr ? mem_857 : _GEN_856; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_858 = 10'h35a == io_addr ? mem_858 : _GEN_857; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_859 = 10'h35b == io_addr ? mem_859 : _GEN_858; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_860 = 10'h35c == io_addr ? mem_860 : _GEN_859; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_861 = 10'h35d == io_addr ? mem_861 : _GEN_860; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_862 = 10'h35e == io_addr ? mem_862 : _GEN_861; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_863 = 10'h35f == io_addr ? mem_863 : _GEN_862; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_864 = 10'h360 == io_addr ? mem_864 : _GEN_863; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_865 = 10'h361 == io_addr ? mem_865 : _GEN_864; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_866 = 10'h362 == io_addr ? mem_866 : _GEN_865; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_867 = 10'h363 == io_addr ? mem_867 : _GEN_866; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_868 = 10'h364 == io_addr ? mem_868 : _GEN_867; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_869 = 10'h365 == io_addr ? mem_869 : _GEN_868; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_870 = 10'h366 == io_addr ? mem_870 : _GEN_869; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_871 = 10'h367 == io_addr ? mem_871 : _GEN_870; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_872 = 10'h368 == io_addr ? mem_872 : _GEN_871; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_873 = 10'h369 == io_addr ? mem_873 : _GEN_872; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_874 = 10'h36a == io_addr ? mem_874 : _GEN_873; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_875 = 10'h36b == io_addr ? mem_875 : _GEN_874; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_876 = 10'h36c == io_addr ? mem_876 : _GEN_875; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_877 = 10'h36d == io_addr ? mem_877 : _GEN_876; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_878 = 10'h36e == io_addr ? mem_878 : _GEN_877; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_879 = 10'h36f == io_addr ? mem_879 : _GEN_878; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_880 = 10'h370 == io_addr ? mem_880 : _GEN_879; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_881 = 10'h371 == io_addr ? mem_881 : _GEN_880; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_882 = 10'h372 == io_addr ? mem_882 : _GEN_881; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_883 = 10'h373 == io_addr ? mem_883 : _GEN_882; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_884 = 10'h374 == io_addr ? mem_884 : _GEN_883; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_885 = 10'h375 == io_addr ? mem_885 : _GEN_884; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_886 = 10'h376 == io_addr ? mem_886 : _GEN_885; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_887 = 10'h377 == io_addr ? mem_887 : _GEN_886; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_888 = 10'h378 == io_addr ? mem_888 : _GEN_887; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_889 = 10'h379 == io_addr ? mem_889 : _GEN_888; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_890 = 10'h37a == io_addr ? mem_890 : _GEN_889; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_891 = 10'h37b == io_addr ? mem_891 : _GEN_890; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_892 = 10'h37c == io_addr ? mem_892 : _GEN_891; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_893 = 10'h37d == io_addr ? mem_893 : _GEN_892; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_894 = 10'h37e == io_addr ? mem_894 : _GEN_893; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_895 = 10'h37f == io_addr ? mem_895 : _GEN_894; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_896 = 10'h380 == io_addr ? mem_896 : _GEN_895; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_897 = 10'h381 == io_addr ? mem_897 : _GEN_896; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_898 = 10'h382 == io_addr ? mem_898 : _GEN_897; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_899 = 10'h383 == io_addr ? mem_899 : _GEN_898; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_900 = 10'h384 == io_addr ? mem_900 : _GEN_899; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_901 = 10'h385 == io_addr ? mem_901 : _GEN_900; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_902 = 10'h386 == io_addr ? mem_902 : _GEN_901; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_903 = 10'h387 == io_addr ? mem_903 : _GEN_902; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_904 = 10'h388 == io_addr ? mem_904 : _GEN_903; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_905 = 10'h389 == io_addr ? mem_905 : _GEN_904; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_906 = 10'h38a == io_addr ? mem_906 : _GEN_905; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_907 = 10'h38b == io_addr ? mem_907 : _GEN_906; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_908 = 10'h38c == io_addr ? mem_908 : _GEN_907; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_909 = 10'h38d == io_addr ? mem_909 : _GEN_908; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_910 = 10'h38e == io_addr ? mem_910 : _GEN_909; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_911 = 10'h38f == io_addr ? mem_911 : _GEN_910; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_912 = 10'h390 == io_addr ? mem_912 : _GEN_911; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_913 = 10'h391 == io_addr ? mem_913 : _GEN_912; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_914 = 10'h392 == io_addr ? mem_914 : _GEN_913; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_915 = 10'h393 == io_addr ? mem_915 : _GEN_914; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_916 = 10'h394 == io_addr ? mem_916 : _GEN_915; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_917 = 10'h395 == io_addr ? mem_917 : _GEN_916; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_918 = 10'h396 == io_addr ? mem_918 : _GEN_917; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_919 = 10'h397 == io_addr ? mem_919 : _GEN_918; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_920 = 10'h398 == io_addr ? mem_920 : _GEN_919; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_921 = 10'h399 == io_addr ? mem_921 : _GEN_920; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_922 = 10'h39a == io_addr ? mem_922 : _GEN_921; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_923 = 10'h39b == io_addr ? mem_923 : _GEN_922; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_924 = 10'h39c == io_addr ? mem_924 : _GEN_923; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_925 = 10'h39d == io_addr ? mem_925 : _GEN_924; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_926 = 10'h39e == io_addr ? mem_926 : _GEN_925; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_927 = 10'h39f == io_addr ? mem_927 : _GEN_926; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_928 = 10'h3a0 == io_addr ? mem_928 : _GEN_927; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_929 = 10'h3a1 == io_addr ? mem_929 : _GEN_928; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_930 = 10'h3a2 == io_addr ? mem_930 : _GEN_929; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_931 = 10'h3a3 == io_addr ? mem_931 : _GEN_930; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_932 = 10'h3a4 == io_addr ? mem_932 : _GEN_931; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_933 = 10'h3a5 == io_addr ? mem_933 : _GEN_932; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_934 = 10'h3a6 == io_addr ? mem_934 : _GEN_933; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_935 = 10'h3a7 == io_addr ? mem_935 : _GEN_934; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_936 = 10'h3a8 == io_addr ? mem_936 : _GEN_935; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_937 = 10'h3a9 == io_addr ? mem_937 : _GEN_936; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_938 = 10'h3aa == io_addr ? mem_938 : _GEN_937; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_939 = 10'h3ab == io_addr ? mem_939 : _GEN_938; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_940 = 10'h3ac == io_addr ? mem_940 : _GEN_939; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_941 = 10'h3ad == io_addr ? mem_941 : _GEN_940; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_942 = 10'h3ae == io_addr ? mem_942 : _GEN_941; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_943 = 10'h3af == io_addr ? mem_943 : _GEN_942; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_944 = 10'h3b0 == io_addr ? mem_944 : _GEN_943; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_945 = 10'h3b1 == io_addr ? mem_945 : _GEN_944; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_946 = 10'h3b2 == io_addr ? mem_946 : _GEN_945; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_947 = 10'h3b3 == io_addr ? mem_947 : _GEN_946; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_948 = 10'h3b4 == io_addr ? mem_948 : _GEN_947; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_949 = 10'h3b5 == io_addr ? mem_949 : _GEN_948; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_950 = 10'h3b6 == io_addr ? mem_950 : _GEN_949; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_951 = 10'h3b7 == io_addr ? mem_951 : _GEN_950; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_952 = 10'h3b8 == io_addr ? mem_952 : _GEN_951; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_953 = 10'h3b9 == io_addr ? mem_953 : _GEN_952; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_954 = 10'h3ba == io_addr ? mem_954 : _GEN_953; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_955 = 10'h3bb == io_addr ? mem_955 : _GEN_954; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_956 = 10'h3bc == io_addr ? mem_956 : _GEN_955; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_957 = 10'h3bd == io_addr ? mem_957 : _GEN_956; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_958 = 10'h3be == io_addr ? mem_958 : _GEN_957; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_959 = 10'h3bf == io_addr ? mem_959 : _GEN_958; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_960 = 10'h3c0 == io_addr ? mem_960 : _GEN_959; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_961 = 10'h3c1 == io_addr ? mem_961 : _GEN_960; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_962 = 10'h3c2 == io_addr ? mem_962 : _GEN_961; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_963 = 10'h3c3 == io_addr ? mem_963 : _GEN_962; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_964 = 10'h3c4 == io_addr ? mem_964 : _GEN_963; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_965 = 10'h3c5 == io_addr ? mem_965 : _GEN_964; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_966 = 10'h3c6 == io_addr ? mem_966 : _GEN_965; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_967 = 10'h3c7 == io_addr ? mem_967 : _GEN_966; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_968 = 10'h3c8 == io_addr ? mem_968 : _GEN_967; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_969 = 10'h3c9 == io_addr ? mem_969 : _GEN_968; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_970 = 10'h3ca == io_addr ? mem_970 : _GEN_969; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_971 = 10'h3cb == io_addr ? mem_971 : _GEN_970; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_972 = 10'h3cc == io_addr ? mem_972 : _GEN_971; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_973 = 10'h3cd == io_addr ? mem_973 : _GEN_972; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_974 = 10'h3ce == io_addr ? mem_974 : _GEN_973; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_975 = 10'h3cf == io_addr ? mem_975 : _GEN_974; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_976 = 10'h3d0 == io_addr ? mem_976 : _GEN_975; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_977 = 10'h3d1 == io_addr ? mem_977 : _GEN_976; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_978 = 10'h3d2 == io_addr ? mem_978 : _GEN_977; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_979 = 10'h3d3 == io_addr ? mem_979 : _GEN_978; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_980 = 10'h3d4 == io_addr ? mem_980 : _GEN_979; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_981 = 10'h3d5 == io_addr ? mem_981 : _GEN_980; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_982 = 10'h3d6 == io_addr ? mem_982 : _GEN_981; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_983 = 10'h3d7 == io_addr ? mem_983 : _GEN_982; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_984 = 10'h3d8 == io_addr ? mem_984 : _GEN_983; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_985 = 10'h3d9 == io_addr ? mem_985 : _GEN_984; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_986 = 10'h3da == io_addr ? mem_986 : _GEN_985; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_987 = 10'h3db == io_addr ? mem_987 : _GEN_986; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_988 = 10'h3dc == io_addr ? mem_988 : _GEN_987; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_989 = 10'h3dd == io_addr ? mem_989 : _GEN_988; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_990 = 10'h3de == io_addr ? mem_990 : _GEN_989; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_991 = 10'h3df == io_addr ? mem_991 : _GEN_990; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_992 = 10'h3e0 == io_addr ? mem_992 : _GEN_991; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_993 = 10'h3e1 == io_addr ? mem_993 : _GEN_992; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_994 = 10'h3e2 == io_addr ? mem_994 : _GEN_993; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_995 = 10'h3e3 == io_addr ? mem_995 : _GEN_994; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_996 = 10'h3e4 == io_addr ? mem_996 : _GEN_995; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_997 = 10'h3e5 == io_addr ? mem_997 : _GEN_996; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_998 = 10'h3e6 == io_addr ? mem_998 : _GEN_997; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_999 = 10'h3e7 == io_addr ? mem_999 : _GEN_998; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1000 = 10'h3e8 == io_addr ? mem_1000 : _GEN_999; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1001 = 10'h3e9 == io_addr ? mem_1001 : _GEN_1000; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1002 = 10'h3ea == io_addr ? mem_1002 : _GEN_1001; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1003 = 10'h3eb == io_addr ? mem_1003 : _GEN_1002; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1004 = 10'h3ec == io_addr ? mem_1004 : _GEN_1003; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1005 = 10'h3ed == io_addr ? mem_1005 : _GEN_1004; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1006 = 10'h3ee == io_addr ? mem_1006 : _GEN_1005; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1007 = 10'h3ef == io_addr ? mem_1007 : _GEN_1006; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1008 = 10'h3f0 == io_addr ? mem_1008 : _GEN_1007; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1009 = 10'h3f1 == io_addr ? mem_1009 : _GEN_1008; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1010 = 10'h3f2 == io_addr ? mem_1010 : _GEN_1009; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1011 = 10'h3f3 == io_addr ? mem_1011 : _GEN_1010; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1012 = 10'h3f4 == io_addr ? mem_1012 : _GEN_1011; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1013 = 10'h3f5 == io_addr ? mem_1013 : _GEN_1012; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1014 = 10'h3f6 == io_addr ? mem_1014 : _GEN_1013; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1015 = 10'h3f7 == io_addr ? mem_1015 : _GEN_1014; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1016 = 10'h3f8 == io_addr ? mem_1016 : _GEN_1015; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1017 = 10'h3f9 == io_addr ? mem_1017 : _GEN_1016; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1018 = 10'h3fa == io_addr ? mem_1018 : _GEN_1017; // @[DataMemoryTest.scala 19:{24,24}]
  wire [31:0] _GEN_1019 = 10'h3fb == io_addr ? mem_1019 : _GEN_1018; // @[DataMemoryTest.scala 19:{24,24}]
  reg [31:0] io_dataOut_REG_1; // @[DataMemoryTest.scala 24:26]
  assign io_dataOut = io_enableWrite ? io_dataOut_REG_1 : io_dataOut_REG; // @[DataMemoryTest.scala 19:14 22:23 24:16]
  always @(posedge clock) begin
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_0 <= 32'h0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_0 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1 <= 32'h1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_2 <= 32'h2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_2 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_3 <= 32'h3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_3 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_4 <= 32'h4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_4 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_5 <= 32'h5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_5 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_6 <= 32'h6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_6 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_7 <= 32'h7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_7 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_8 <= 32'h8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_8 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_9 <= 32'h9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_9 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_10 <= 32'ha; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_10 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_11 <= 32'hb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_11 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_12 <= 32'hc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_12 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_13 <= 32'hd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_13 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_14 <= 32'he; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_14 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_15 <= 32'hf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_15 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_16 <= 32'h10; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_16 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_17 <= 32'h11; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_17 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_18 <= 32'h12; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_18 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_19 <= 32'h13; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_19 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_20 <= 32'h14; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_20 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_21 <= 32'h15; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_21 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_22 <= 32'h16; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_22 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_23 <= 32'h17; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_23 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_24 <= 32'h18; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_24 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_25 <= 32'h19; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_25 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_26 <= 32'h1a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_26 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_27 <= 32'h1b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_27 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_28 <= 32'h1c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_28 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_29 <= 32'h1d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_29 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_30 <= 32'h1e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_30 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_31 <= 32'h1f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_31 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_32 <= 32'h20; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_32 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_33 <= 32'h21; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_33 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_34 <= 32'h22; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_34 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_35 <= 32'h23; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_35 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_36 <= 32'h24; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_36 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_37 <= 32'h25; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_37 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_38 <= 32'h26; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_38 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_39 <= 32'h27; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_39 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_40 <= 32'h28; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_40 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_41 <= 32'h29; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_41 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_42 <= 32'h2a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_42 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_43 <= 32'h2b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_43 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_44 <= 32'h2c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_44 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_45 <= 32'h2d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_45 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_46 <= 32'h2e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_46 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_47 <= 32'h2f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_47 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_48 <= 32'h30; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_48 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_49 <= 32'h31; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_49 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_50 <= 32'h32; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_50 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_51 <= 32'h33; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_51 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_52 <= 32'h34; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_52 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_53 <= 32'h35; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_53 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_54 <= 32'h36; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_54 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_55 <= 32'h37; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_55 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_56 <= 32'h38; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_56 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_57 <= 32'h39; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_57 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_58 <= 32'h3a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_58 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_59 <= 32'h3b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_59 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_60 <= 32'h3c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_60 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_61 <= 32'h3d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_61 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_62 <= 32'h3e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_62 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_63 <= 32'h3f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_63 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_64 <= 32'h40; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h40 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_64 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_65 <= 32'h41; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h41 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_65 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_66 <= 32'h42; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h42 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_66 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_67 <= 32'h43; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h43 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_67 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_68 <= 32'h44; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h44 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_68 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_69 <= 32'h45; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h45 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_69 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_70 <= 32'h46; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h46 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_70 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_71 <= 32'h47; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h47 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_71 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_72 <= 32'h48; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h48 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_72 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_73 <= 32'h49; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h49 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_73 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_74 <= 32'h4a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_74 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_75 <= 32'h4b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_75 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_76 <= 32'h4c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_76 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_77 <= 32'h4d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_77 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_78 <= 32'h4e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_78 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_79 <= 32'h4f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h4f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_79 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_80 <= 32'h50; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h50 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_80 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_81 <= 32'h51; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h51 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_81 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_82 <= 32'h52; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h52 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_82 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_83 <= 32'h53; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h53 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_83 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_84 <= 32'h54; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h54 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_84 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_85 <= 32'h55; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h55 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_85 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_86 <= 32'h56; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h56 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_86 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_87 <= 32'h57; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h57 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_87 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_88 <= 32'h58; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h58 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_88 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_89 <= 32'h59; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h59 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_89 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_90 <= 32'h5a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_90 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_91 <= 32'h5b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_91 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_92 <= 32'h5c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_92 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_93 <= 32'h5d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_93 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_94 <= 32'h5e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_94 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_95 <= 32'h5f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h5f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_95 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_96 <= 32'h60; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h60 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_96 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_97 <= 32'h61; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h61 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_97 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_98 <= 32'h62; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h62 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_98 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_99 <= 32'h63; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h63 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_99 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_100 <= 32'h64; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h64 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_100 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_101 <= 32'h65; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h65 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_101 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_102 <= 32'h66; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h66 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_102 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_103 <= 32'h67; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h67 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_103 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_104 <= 32'h68; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h68 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_104 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_105 <= 32'h69; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h69 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_105 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_106 <= 32'h6a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_106 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_107 <= 32'h6b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_107 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_108 <= 32'h6c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_108 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_109 <= 32'h6d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_109 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_110 <= 32'h6e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_110 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_111 <= 32'h6f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h6f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_111 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_112 <= 32'h70; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h70 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_112 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_113 <= 32'h71; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h71 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_113 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_114 <= 32'h72; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h72 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_114 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_115 <= 32'h73; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h73 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_115 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_116 <= 32'h74; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h74 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_116 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_117 <= 32'h75; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h75 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_117 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_118 <= 32'h76; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h76 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_118 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_119 <= 32'h77; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h77 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_119 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_120 <= 32'h78; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h78 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_120 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_121 <= 32'h79; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h79 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_121 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_122 <= 32'h7a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_122 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_123 <= 32'h7b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_123 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_124 <= 32'h7c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_124 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_125 <= 32'h7d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_125 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_126 <= 32'h7e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_126 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_127 <= 32'h7f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h7f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_127 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_128 <= 32'h80; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h80 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_128 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_129 <= 32'h81; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h81 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_129 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_130 <= 32'h82; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h82 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_130 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_131 <= 32'h83; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h83 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_131 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_132 <= 32'h84; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h84 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_132 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_133 <= 32'h85; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h85 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_133 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_134 <= 32'h86; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h86 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_134 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_135 <= 32'h87; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h87 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_135 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_136 <= 32'h88; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h88 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_136 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_137 <= 32'h89; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h89 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_137 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_138 <= 32'h8a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_138 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_139 <= 32'h8b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_139 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_140 <= 32'h8c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_140 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_141 <= 32'h8d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_141 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_142 <= 32'h8e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_142 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_143 <= 32'h8f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h8f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_143 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_144 <= 32'h90; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h90 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_144 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_145 <= 32'h91; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h91 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_145 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_146 <= 32'h92; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h92 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_146 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_147 <= 32'h93; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h93 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_147 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_148 <= 32'h94; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h94 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_148 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_149 <= 32'h95; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h95 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_149 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_150 <= 32'h96; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h96 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_150 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_151 <= 32'h97; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h97 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_151 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_152 <= 32'h98; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h98 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_152 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_153 <= 32'h99; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h99 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_153 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_154 <= 32'h9a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_154 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_155 <= 32'h9b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_155 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_156 <= 32'h9c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_156 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_157 <= 32'h9d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_157 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_158 <= 32'h9e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_158 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_159 <= 32'h9f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h9f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_159 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_160 <= 32'ha0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_160 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_161 <= 32'ha1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_161 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_162 <= 32'ha2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_162 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_163 <= 32'ha3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_163 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_164 <= 32'ha4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_164 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_165 <= 32'ha5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_165 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_166 <= 32'ha6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_166 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_167 <= 32'ha7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_167 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_168 <= 32'ha8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_168 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_169 <= 32'ha9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'ha9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_169 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_170 <= 32'haa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'haa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_170 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_171 <= 32'hab; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hab == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_171 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_172 <= 32'hac; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hac == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_172 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_173 <= 32'had; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'had == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_173 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_174 <= 32'hae; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hae == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_174 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_175 <= 32'haf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'haf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_175 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_176 <= 32'hb0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_176 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_177 <= 32'hb1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_177 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_178 <= 32'hb2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_178 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_179 <= 32'hb3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_179 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_180 <= 32'hb4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_180 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_181 <= 32'hb5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_181 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_182 <= 32'hb6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_182 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_183 <= 32'hb7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_183 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_184 <= 32'hb8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_184 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_185 <= 32'hb9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hb9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_185 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_186 <= 32'hba; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hba == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_186 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_187 <= 32'hbb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hbb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_187 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_188 <= 32'hbc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hbc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_188 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_189 <= 32'hbd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hbd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_189 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_190 <= 32'hbe; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hbe == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_190 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_191 <= 32'hbf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hbf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_191 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_192 <= 32'hc0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_192 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_193 <= 32'hc1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_193 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_194 <= 32'hc2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_194 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_195 <= 32'hc3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_195 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_196 <= 32'hc4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_196 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_197 <= 32'hc5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_197 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_198 <= 32'hc6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_198 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_199 <= 32'hc7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_199 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_200 <= 32'hc8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_200 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_201 <= 32'hc9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hc9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_201 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_202 <= 32'hca; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hca == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_202 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_203 <= 32'hcb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hcb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_203 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_204 <= 32'hcc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hcc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_204 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_205 <= 32'hcd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hcd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_205 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_206 <= 32'hce; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hce == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_206 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_207 <= 32'hcf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hcf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_207 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_208 <= 32'hd0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_208 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_209 <= 32'hd1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_209 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_210 <= 32'hd2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_210 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_211 <= 32'hd3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_211 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_212 <= 32'hd4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_212 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_213 <= 32'hd5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_213 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_214 <= 32'hd6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_214 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_215 <= 32'hd7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_215 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_216 <= 32'hd8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_216 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_217 <= 32'hd9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hd9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_217 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_218 <= 32'hda; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hda == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_218 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_219 <= 32'hdb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hdb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_219 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_220 <= 32'hdc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hdc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_220 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_221 <= 32'hdd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hdd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_221 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_222 <= 32'hde; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hde == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_222 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_223 <= 32'hdf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hdf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_223 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_224 <= 32'he0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_224 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_225 <= 32'he1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_225 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_226 <= 32'he2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_226 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_227 <= 32'he3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_227 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_228 <= 32'he4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_228 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_229 <= 32'he5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_229 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_230 <= 32'he6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_230 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_231 <= 32'he7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_231 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_232 <= 32'he8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_232 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_233 <= 32'he9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'he9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_233 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_234 <= 32'hea; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hea == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_234 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_235 <= 32'heb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'heb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_235 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_236 <= 32'hec; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hec == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_236 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_237 <= 32'hed; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hed == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_237 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_238 <= 32'hee; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hee == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_238 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_239 <= 32'hef; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hef == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_239 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_240 <= 32'hf0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_240 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_241 <= 32'hf1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_241 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_242 <= 32'hf2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_242 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_243 <= 32'hf3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_243 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_244 <= 32'hf4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_244 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_245 <= 32'hf5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_245 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_246 <= 32'hf6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_246 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_247 <= 32'hf7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_247 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_248 <= 32'hf8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_248 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_249 <= 32'hf9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hf9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_249 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_250 <= 32'hfa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hfa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_250 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_251 <= 32'hfb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hfb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_251 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_252 <= 32'hfc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hfc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_252 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_253 <= 32'hfd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hfd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_253 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_254 <= 32'hfe; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hfe == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_254 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_255 <= 32'hff; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'hff == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_255 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_256 <= 32'h100; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h100 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_256 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_257 <= 32'h101; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h101 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_257 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_258 <= 32'h102; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h102 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_258 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_259 <= 32'h103; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h103 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_259 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_260 <= 32'h104; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h104 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_260 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_261 <= 32'h105; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h105 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_261 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_262 <= 32'h106; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h106 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_262 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_263 <= 32'h107; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h107 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_263 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_264 <= 32'h108; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h108 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_264 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_265 <= 32'h109; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h109 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_265 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_266 <= 32'h10a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_266 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_267 <= 32'h10b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_267 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_268 <= 32'h10c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_268 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_269 <= 32'h10d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_269 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_270 <= 32'h10e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_270 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_271 <= 32'h10f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h10f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_271 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_272 <= 32'h110; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h110 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_272 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_273 <= 32'h111; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h111 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_273 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_274 <= 32'h112; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h112 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_274 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_275 <= 32'h113; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h113 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_275 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_276 <= 32'h114; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h114 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_276 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_277 <= 32'h115; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h115 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_277 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_278 <= 32'h116; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h116 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_278 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_279 <= 32'h117; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h117 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_279 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_280 <= 32'h118; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h118 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_280 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_281 <= 32'h119; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h119 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_281 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_282 <= 32'h11a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_282 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_283 <= 32'h11b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_283 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_284 <= 32'h11c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_284 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_285 <= 32'h11d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_285 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_286 <= 32'h11e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_286 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_287 <= 32'h11f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h11f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_287 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_288 <= 32'h120; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h120 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_288 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_289 <= 32'h121; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h121 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_289 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_290 <= 32'h122; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h122 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_290 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_291 <= 32'h123; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h123 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_291 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_292 <= 32'h124; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h124 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_292 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_293 <= 32'h125; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h125 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_293 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_294 <= 32'h126; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h126 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_294 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_295 <= 32'h127; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h127 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_295 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_296 <= 32'h128; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h128 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_296 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_297 <= 32'h129; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h129 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_297 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_298 <= 32'h12a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_298 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_299 <= 32'h12b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_299 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_300 <= 32'h12c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_300 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_301 <= 32'h12d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_301 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_302 <= 32'h12e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_302 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_303 <= 32'h12f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h12f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_303 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_304 <= 32'h130; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h130 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_304 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_305 <= 32'h131; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h131 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_305 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_306 <= 32'h132; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h132 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_306 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_307 <= 32'h133; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h133 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_307 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_308 <= 32'h134; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h134 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_308 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_309 <= 32'h135; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h135 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_309 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_310 <= 32'h136; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h136 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_310 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_311 <= 32'h137; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h137 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_311 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_312 <= 32'h138; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h138 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_312 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_313 <= 32'h139; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h139 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_313 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_314 <= 32'h13a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_314 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_315 <= 32'h13b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_315 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_316 <= 32'h13c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_316 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_317 <= 32'h13d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_317 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_318 <= 32'h13e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_318 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_319 <= 32'h13f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h13f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_319 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_320 <= 32'h140; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h140 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_320 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_321 <= 32'h141; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h141 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_321 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_322 <= 32'h142; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h142 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_322 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_323 <= 32'h143; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h143 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_323 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_324 <= 32'h144; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h144 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_324 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_325 <= 32'h145; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h145 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_325 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_326 <= 32'h146; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h146 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_326 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_327 <= 32'h147; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h147 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_327 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_328 <= 32'h148; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h148 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_328 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_329 <= 32'h149; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h149 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_329 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_330 <= 32'h14a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_330 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_331 <= 32'h14b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_331 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_332 <= 32'h14c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_332 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_333 <= 32'h14d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_333 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_334 <= 32'h14e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_334 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_335 <= 32'h14f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h14f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_335 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_336 <= 32'h150; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h150 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_336 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_337 <= 32'h151; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h151 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_337 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_338 <= 32'h152; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h152 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_338 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_339 <= 32'h153; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h153 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_339 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_340 <= 32'h154; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h154 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_340 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_341 <= 32'h155; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h155 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_341 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_342 <= 32'h156; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h156 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_342 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_343 <= 32'h157; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h157 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_343 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_344 <= 32'h158; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h158 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_344 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_345 <= 32'h159; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h159 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_345 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_346 <= 32'h15a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_346 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_347 <= 32'h15b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_347 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_348 <= 32'h15c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_348 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_349 <= 32'h15d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_349 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_350 <= 32'h15e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_350 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_351 <= 32'h15f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h15f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_351 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_352 <= 32'h160; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h160 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_352 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_353 <= 32'h161; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h161 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_353 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_354 <= 32'h162; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h162 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_354 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_355 <= 32'h163; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h163 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_355 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_356 <= 32'h164; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h164 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_356 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_357 <= 32'h165; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h165 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_357 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_358 <= 32'h166; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h166 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_358 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_359 <= 32'h167; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h167 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_359 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_360 <= 32'h168; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h168 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_360 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_361 <= 32'h169; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h169 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_361 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_362 <= 32'h16a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_362 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_363 <= 32'h16b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_363 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_364 <= 32'h16c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_364 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_365 <= 32'h16d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_365 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_366 <= 32'h16e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_366 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_367 <= 32'h16f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h16f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_367 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_368 <= 32'h170; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h170 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_368 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_369 <= 32'h171; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h171 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_369 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_370 <= 32'h172; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h172 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_370 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_371 <= 32'h173; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h173 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_371 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_372 <= 32'h174; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h174 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_372 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_373 <= 32'h175; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h175 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_373 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_374 <= 32'h176; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h176 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_374 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_375 <= 32'h177; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h177 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_375 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_376 <= 32'h178; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h178 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_376 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_377 <= 32'h179; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h179 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_377 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_378 <= 32'h17a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_378 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_379 <= 32'h17b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_379 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_380 <= 32'h17c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_380 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_381 <= 32'h17d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_381 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_382 <= 32'h17e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_382 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_383 <= 32'h17f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h17f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_383 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_384 <= 32'h180; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h180 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_384 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_385 <= 32'h181; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h181 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_385 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_386 <= 32'h182; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h182 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_386 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_387 <= 32'h183; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h183 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_387 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_388 <= 32'h184; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h184 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_388 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_389 <= 32'h185; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h185 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_389 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_390 <= 32'h186; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h186 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_390 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_391 <= 32'h187; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h187 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_391 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_392 <= 32'h188; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h188 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_392 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_393 <= 32'h189; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h189 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_393 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_394 <= 32'h18a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_394 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_395 <= 32'h18b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_395 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_396 <= 32'h18c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_396 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_397 <= 32'h18d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_397 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_398 <= 32'h18e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_398 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_399 <= 32'h18f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h18f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_399 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_400 <= 32'h190; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h190 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_400 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_401 <= 32'h191; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h191 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_401 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_402 <= 32'h192; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h192 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_402 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_403 <= 32'h193; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h193 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_403 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_404 <= 32'h194; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h194 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_404 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_405 <= 32'h195; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h195 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_405 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_406 <= 32'h196; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h196 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_406 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_407 <= 32'h197; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h197 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_407 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_408 <= 32'h198; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h198 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_408 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_409 <= 32'h199; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h199 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_409 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_410 <= 32'h19a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_410 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_411 <= 32'h19b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_411 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_412 <= 32'h19c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_412 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_413 <= 32'h19d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_413 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_414 <= 32'h19e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_414 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_415 <= 32'h19f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h19f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_415 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_416 <= 32'h1a0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_416 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_417 <= 32'h1a1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_417 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_418 <= 32'h1a2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_418 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_419 <= 32'h1a3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_419 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_420 <= 32'h1a4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_420 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_421 <= 32'h1a5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_421 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_422 <= 32'h1a6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_422 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_423 <= 32'h1a7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_423 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_424 <= 32'h1a8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_424 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_425 <= 32'h1a9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1a9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_425 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_426 <= 32'h1aa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1aa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_426 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_427 <= 32'h1ab; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ab == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_427 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_428 <= 32'h1ac; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ac == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_428 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_429 <= 32'h1ad; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ad == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_429 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_430 <= 32'h1ae; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ae == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_430 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_431 <= 32'h1af; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1af == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_431 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_432 <= 32'h1b0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_432 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_433 <= 32'h1b1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_433 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_434 <= 32'h1b2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_434 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_435 <= 32'h1b3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_435 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_436 <= 32'h1b4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_436 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_437 <= 32'h1b5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_437 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_438 <= 32'h1b6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_438 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_439 <= 32'h1b7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_439 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_440 <= 32'h1b8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_440 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_441 <= 32'h1b9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1b9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_441 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_442 <= 32'h1ba; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ba == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_442 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_443 <= 32'h1bb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1bb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_443 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_444 <= 32'h1bc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1bc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_444 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_445 <= 32'h1bd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1bd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_445 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_446 <= 32'h1be; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1be == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_446 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_447 <= 32'h1bf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1bf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_447 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_448 <= 32'h1c0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_448 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_449 <= 32'h1c1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_449 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_450 <= 32'h1c2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_450 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_451 <= 32'h1c3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_451 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_452 <= 32'h1c4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_452 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_453 <= 32'h1c5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_453 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_454 <= 32'h1c6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_454 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_455 <= 32'h1c7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_455 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_456 <= 32'h1c8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_456 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_457 <= 32'h1c9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1c9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_457 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_458 <= 32'h1ca; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ca == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_458 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_459 <= 32'h1cb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1cb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_459 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_460 <= 32'h1cc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1cc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_460 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_461 <= 32'h1cd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1cd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_461 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_462 <= 32'h1ce; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ce == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_462 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_463 <= 32'h1cf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1cf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_463 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_464 <= 32'h1d0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_464 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_465 <= 32'h1d1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_465 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_466 <= 32'h1d2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_466 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_467 <= 32'h1d3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_467 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_468 <= 32'h1d4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_468 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_469 <= 32'h1d5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_469 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_470 <= 32'h1d6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_470 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_471 <= 32'h1d7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_471 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_472 <= 32'h1d8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_472 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_473 <= 32'h1d9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1d9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_473 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_474 <= 32'h1da; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1da == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_474 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_475 <= 32'h1db; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1db == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_475 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_476 <= 32'h1dc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1dc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_476 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_477 <= 32'h1dd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1dd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_477 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_478 <= 32'h1de; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1de == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_478 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_479 <= 32'h1df; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1df == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_479 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_480 <= 32'h1e0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_480 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_481 <= 32'h1e1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_481 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_482 <= 32'h1e2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_482 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_483 <= 32'h1e3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_483 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_484 <= 32'h1e4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_484 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_485 <= 32'h1e5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_485 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_486 <= 32'h1e6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_486 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_487 <= 32'h1e7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_487 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_488 <= 32'h1e8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_488 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_489 <= 32'h1e9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1e9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_489 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_490 <= 32'h1ea; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ea == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_490 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_491 <= 32'h1eb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1eb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_491 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_492 <= 32'h1ec; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ec == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_492 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_493 <= 32'h1ed; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ed == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_493 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_494 <= 32'h1ee; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ee == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_494 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_495 <= 32'h1ef; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ef == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_495 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_496 <= 32'h1f0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_496 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_497 <= 32'h1f1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_497 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_498 <= 32'h1f2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_498 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_499 <= 32'h1f3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_499 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_500 <= 32'h1f4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_500 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_501 <= 32'h1f5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_501 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_502 <= 32'h1f6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_502 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_503 <= 32'h1f7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_503 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_504 <= 32'h1f8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_504 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_505 <= 32'h1f9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1f9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_505 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_506 <= 32'h1fa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1fa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_506 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_507 <= 32'h1fb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1fb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_507 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_508 <= 32'h1fc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1fc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_508 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_509 <= 32'h1fd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1fd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_509 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_510 <= 32'h1fe; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1fe == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_510 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_511 <= 32'h1ff; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h1ff == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_511 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_512 <= 32'h200; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h200 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_512 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_513 <= 32'h201; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h201 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_513 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_514 <= 32'h202; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h202 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_514 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_515 <= 32'h203; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h203 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_515 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_516 <= 32'h204; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h204 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_516 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_517 <= 32'h205; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h205 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_517 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_518 <= 32'h206; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h206 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_518 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_519 <= 32'h207; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h207 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_519 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_520 <= 32'h208; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h208 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_520 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_521 <= 32'h209; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h209 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_521 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_522 <= 32'h20a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_522 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_523 <= 32'h20b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_523 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_524 <= 32'h20c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_524 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_525 <= 32'h20d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_525 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_526 <= 32'h20e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_526 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_527 <= 32'h20f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h20f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_527 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_528 <= 32'h210; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h210 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_528 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_529 <= 32'h211; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h211 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_529 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_530 <= 32'h212; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h212 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_530 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_531 <= 32'h213; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h213 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_531 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_532 <= 32'h214; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h214 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_532 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_533 <= 32'h215; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h215 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_533 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_534 <= 32'h216; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h216 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_534 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_535 <= 32'h217; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h217 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_535 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_536 <= 32'h218; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h218 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_536 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_537 <= 32'h219; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h219 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_537 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_538 <= 32'h21a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_538 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_539 <= 32'h21b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_539 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_540 <= 32'h21c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_540 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_541 <= 32'h21d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_541 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_542 <= 32'h21e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_542 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_543 <= 32'h21f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h21f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_543 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_544 <= 32'h220; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h220 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_544 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_545 <= 32'h221; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h221 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_545 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_546 <= 32'h222; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h222 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_546 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_547 <= 32'h223; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h223 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_547 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_548 <= 32'h224; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h224 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_548 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_549 <= 32'h225; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h225 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_549 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_550 <= 32'h226; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h226 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_550 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_551 <= 32'h227; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h227 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_551 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_552 <= 32'h228; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h228 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_552 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_553 <= 32'h229; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h229 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_553 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_554 <= 32'h22a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_554 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_555 <= 32'h22b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_555 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_556 <= 32'h22c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_556 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_557 <= 32'h22d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_557 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_558 <= 32'h22e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_558 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_559 <= 32'h22f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h22f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_559 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_560 <= 32'h230; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h230 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_560 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_561 <= 32'h231; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h231 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_561 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_562 <= 32'h232; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h232 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_562 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_563 <= 32'h233; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h233 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_563 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_564 <= 32'h234; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h234 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_564 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_565 <= 32'h235; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h235 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_565 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_566 <= 32'h236; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h236 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_566 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_567 <= 32'h237; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h237 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_567 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_568 <= 32'h238; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h238 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_568 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_569 <= 32'h239; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h239 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_569 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_570 <= 32'h23a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_570 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_571 <= 32'h23b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_571 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_572 <= 32'h23c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_572 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_573 <= 32'h23d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_573 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_574 <= 32'h23e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_574 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_575 <= 32'h23f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h23f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_575 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_576 <= 32'h240; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h240 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_576 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_577 <= 32'h241; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h241 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_577 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_578 <= 32'h242; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h242 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_578 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_579 <= 32'h243; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h243 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_579 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_580 <= 32'h244; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h244 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_580 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_581 <= 32'h245; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h245 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_581 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_582 <= 32'h246; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h246 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_582 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_583 <= 32'h247; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h247 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_583 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_584 <= 32'h248; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h248 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_584 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_585 <= 32'h249; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h249 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_585 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_586 <= 32'h24a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_586 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_587 <= 32'h24b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_587 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_588 <= 32'h24c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_588 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_589 <= 32'h24d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_589 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_590 <= 32'h24e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_590 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_591 <= 32'h24f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h24f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_591 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_592 <= 32'h250; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h250 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_592 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_593 <= 32'h251; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h251 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_593 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_594 <= 32'h252; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h252 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_594 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_595 <= 32'h253; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h253 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_595 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_596 <= 32'h254; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h254 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_596 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_597 <= 32'h255; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h255 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_597 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_598 <= 32'h256; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h256 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_598 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_599 <= 32'h257; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h257 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_599 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_600 <= 32'h258; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h258 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_600 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_601 <= 32'h259; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h259 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_601 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_602 <= 32'h25a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_602 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_603 <= 32'h25b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_603 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_604 <= 32'h25c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_604 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_605 <= 32'h25d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_605 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_606 <= 32'h25e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_606 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_607 <= 32'h25f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h25f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_607 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_608 <= 32'h260; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h260 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_608 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_609 <= 32'h261; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h261 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_609 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_610 <= 32'h262; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h262 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_610 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_611 <= 32'h263; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h263 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_611 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_612 <= 32'h264; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h264 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_612 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_613 <= 32'h265; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h265 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_613 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_614 <= 32'h266; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h266 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_614 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_615 <= 32'h267; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h267 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_615 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_616 <= 32'h268; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h268 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_616 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_617 <= 32'h269; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h269 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_617 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_618 <= 32'h26a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_618 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_619 <= 32'h26b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_619 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_620 <= 32'h26c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_620 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_621 <= 32'h26d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_621 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_622 <= 32'h26e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_622 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_623 <= 32'h26f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h26f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_623 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_624 <= 32'h270; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h270 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_624 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_625 <= 32'h271; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h271 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_625 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_626 <= 32'h272; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h272 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_626 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_627 <= 32'h273; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h273 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_627 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_628 <= 32'h274; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h274 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_628 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_629 <= 32'h275; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h275 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_629 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_630 <= 32'h276; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h276 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_630 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_631 <= 32'h277; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h277 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_631 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_632 <= 32'h278; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h278 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_632 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_633 <= 32'h279; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h279 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_633 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_634 <= 32'h27a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_634 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_635 <= 32'h27b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_635 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_636 <= 32'h27c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_636 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_637 <= 32'h27d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_637 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_638 <= 32'h27e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_638 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_639 <= 32'h27f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h27f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_639 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_640 <= 32'h280; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h280 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_640 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_641 <= 32'h281; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h281 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_641 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_642 <= 32'h282; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h282 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_642 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_643 <= 32'h283; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h283 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_643 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_644 <= 32'h284; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h284 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_644 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_645 <= 32'h285; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h285 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_645 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_646 <= 32'h286; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h286 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_646 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_647 <= 32'h287; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h287 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_647 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_648 <= 32'h288; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h288 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_648 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_649 <= 32'h289; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h289 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_649 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_650 <= 32'h28a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_650 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_651 <= 32'h28b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_651 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_652 <= 32'h28c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_652 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_653 <= 32'h28d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_653 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_654 <= 32'h28e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_654 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_655 <= 32'h28f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h28f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_655 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_656 <= 32'h290; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h290 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_656 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_657 <= 32'h291; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h291 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_657 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_658 <= 32'h292; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h292 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_658 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_659 <= 32'h293; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h293 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_659 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_660 <= 32'h294; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h294 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_660 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_661 <= 32'h295; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h295 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_661 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_662 <= 32'h296; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h296 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_662 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_663 <= 32'h297; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h297 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_663 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_664 <= 32'h298; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h298 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_664 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_665 <= 32'h299; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h299 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_665 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_666 <= 32'h29a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_666 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_667 <= 32'h29b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_667 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_668 <= 32'h29c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_668 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_669 <= 32'h29d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_669 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_670 <= 32'h29e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_670 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_671 <= 32'h29f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h29f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_671 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_672 <= 32'h2a0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_672 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_673 <= 32'h2a1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_673 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_674 <= 32'h2a2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_674 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_675 <= 32'h2a3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_675 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_676 <= 32'h2a4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_676 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_677 <= 32'h2a5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_677 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_678 <= 32'h2a6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_678 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_679 <= 32'h2a7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_679 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_680 <= 32'h2a8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_680 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_681 <= 32'h2a9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2a9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_681 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_682 <= 32'h2aa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2aa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_682 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_683 <= 32'h2ab; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ab == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_683 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_684 <= 32'h2ac; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ac == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_684 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_685 <= 32'h2ad; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ad == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_685 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_686 <= 32'h2ae; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ae == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_686 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_687 <= 32'h2af; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2af == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_687 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_688 <= 32'h2b0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_688 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_689 <= 32'h2b1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_689 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_690 <= 32'h2b2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_690 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_691 <= 32'h2b3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_691 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_692 <= 32'h2b4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_692 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_693 <= 32'h2b5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_693 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_694 <= 32'h2b6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_694 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_695 <= 32'h2b7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_695 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_696 <= 32'h2b8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_696 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_697 <= 32'h2b9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2b9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_697 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_698 <= 32'h2ba; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ba == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_698 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_699 <= 32'h2bb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2bb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_699 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_700 <= 32'h2bc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2bc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_700 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_701 <= 32'h2bd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2bd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_701 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_702 <= 32'h2be; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2be == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_702 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_703 <= 32'h2bf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2bf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_703 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_704 <= 32'h2c0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_704 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_705 <= 32'h2c1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_705 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_706 <= 32'h2c2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_706 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_707 <= 32'h2c3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_707 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_708 <= 32'h2c4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_708 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_709 <= 32'h2c5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_709 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_710 <= 32'h2c6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_710 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_711 <= 32'h2c7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_711 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_712 <= 32'h2c8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_712 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_713 <= 32'h2c9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2c9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_713 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_714 <= 32'h2ca; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ca == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_714 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_715 <= 32'h2cb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2cb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_715 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_716 <= 32'h2cc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2cc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_716 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_717 <= 32'h2cd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2cd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_717 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_718 <= 32'h2ce; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ce == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_718 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_719 <= 32'h2cf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2cf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_719 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_720 <= 32'h2d0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_720 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_721 <= 32'h2d1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_721 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_722 <= 32'h2d2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_722 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_723 <= 32'h2d3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_723 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_724 <= 32'h2d4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_724 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_725 <= 32'h2d5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_725 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_726 <= 32'h2d6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_726 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_727 <= 32'h2d7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_727 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_728 <= 32'h2d8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_728 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_729 <= 32'h2d9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2d9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_729 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_730 <= 32'h2da; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2da == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_730 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_731 <= 32'h2db; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2db == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_731 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_732 <= 32'h2dc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2dc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_732 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_733 <= 32'h2dd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2dd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_733 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_734 <= 32'h2de; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2de == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_734 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_735 <= 32'h2df; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2df == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_735 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_736 <= 32'h2e0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_736 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_737 <= 32'h2e1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_737 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_738 <= 32'h2e2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_738 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_739 <= 32'h2e3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_739 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_740 <= 32'h2e4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_740 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_741 <= 32'h2e5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_741 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_742 <= 32'h2e6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_742 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_743 <= 32'h2e7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_743 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_744 <= 32'h2e8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_744 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_745 <= 32'h2e9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2e9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_745 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_746 <= 32'h2ea; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ea == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_746 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_747 <= 32'h2eb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2eb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_747 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_748 <= 32'h2ec; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ec == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_748 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_749 <= 32'h2ed; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ed == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_749 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_750 <= 32'h2ee; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ee == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_750 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_751 <= 32'h2ef; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ef == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_751 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_752 <= 32'h2f0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_752 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_753 <= 32'h2f1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_753 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_754 <= 32'h2f2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_754 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_755 <= 32'h2f3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_755 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_756 <= 32'h2f4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_756 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_757 <= 32'h2f5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_757 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_758 <= 32'h2f6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_758 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_759 <= 32'h2f7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_759 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_760 <= 32'h2f8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_760 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_761 <= 32'h2f9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2f9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_761 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_762 <= 32'h2fa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2fa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_762 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_763 <= 32'h2fb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2fb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_763 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_764 <= 32'h2fc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2fc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_764 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_765 <= 32'h2fd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2fd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_765 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_766 <= 32'h2fe; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2fe == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_766 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_767 <= 32'h2ff; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h2ff == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_767 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_768 <= 32'h300; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h300 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_768 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_769 <= 32'h301; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h301 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_769 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_770 <= 32'h302; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h302 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_770 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_771 <= 32'h303; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h303 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_771 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_772 <= 32'h304; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h304 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_772 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_773 <= 32'h305; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h305 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_773 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_774 <= 32'h306; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h306 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_774 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_775 <= 32'h307; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h307 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_775 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_776 <= 32'h308; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h308 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_776 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_777 <= 32'h309; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h309 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_777 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_778 <= 32'h30a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_778 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_779 <= 32'h30b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_779 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_780 <= 32'h30c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_780 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_781 <= 32'h30d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_781 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_782 <= 32'h30e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_782 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_783 <= 32'h30f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h30f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_783 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_784 <= 32'h310; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h310 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_784 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_785 <= 32'h311; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h311 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_785 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_786 <= 32'h312; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h312 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_786 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_787 <= 32'h313; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h313 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_787 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_788 <= 32'h314; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h314 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_788 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_789 <= 32'h315; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h315 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_789 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_790 <= 32'h316; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h316 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_790 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_791 <= 32'h317; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h317 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_791 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_792 <= 32'h318; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h318 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_792 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_793 <= 32'h319; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h319 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_793 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_794 <= 32'h31a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_794 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_795 <= 32'h31b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_795 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_796 <= 32'h31c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_796 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_797 <= 32'h31d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_797 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_798 <= 32'h31e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_798 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_799 <= 32'h31f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h31f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_799 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_800 <= 32'h320; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h320 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_800 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_801 <= 32'h321; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h321 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_801 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_802 <= 32'h322; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h322 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_802 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_803 <= 32'h323; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h323 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_803 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_804 <= 32'h324; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h324 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_804 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_805 <= 32'h325; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h325 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_805 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_806 <= 32'h326; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h326 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_806 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_807 <= 32'h327; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h327 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_807 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_808 <= 32'h328; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h328 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_808 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_809 <= 32'h329; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h329 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_809 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_810 <= 32'h32a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_810 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_811 <= 32'h32b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_811 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_812 <= 32'h32c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_812 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_813 <= 32'h32d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_813 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_814 <= 32'h32e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_814 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_815 <= 32'h32f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h32f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_815 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_816 <= 32'h330; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h330 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_816 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_817 <= 32'h331; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h331 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_817 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_818 <= 32'h332; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h332 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_818 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_819 <= 32'h333; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h333 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_819 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_820 <= 32'h334; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h334 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_820 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_821 <= 32'h335; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h335 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_821 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_822 <= 32'h336; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h336 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_822 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_823 <= 32'h337; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h337 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_823 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_824 <= 32'h338; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h338 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_824 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_825 <= 32'h339; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h339 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_825 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_826 <= 32'h33a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_826 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_827 <= 32'h33b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_827 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_828 <= 32'h33c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_828 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_829 <= 32'h33d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_829 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_830 <= 32'h33e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_830 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_831 <= 32'h33f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h33f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_831 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_832 <= 32'h340; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h340 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_832 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_833 <= 32'h341; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h341 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_833 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_834 <= 32'h342; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h342 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_834 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_835 <= 32'h343; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h343 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_835 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_836 <= 32'h344; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h344 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_836 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_837 <= 32'h345; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h345 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_837 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_838 <= 32'h346; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h346 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_838 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_839 <= 32'h347; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h347 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_839 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_840 <= 32'h348; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h348 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_840 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_841 <= 32'h349; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h349 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_841 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_842 <= 32'h34a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_842 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_843 <= 32'h34b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_843 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_844 <= 32'h34c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_844 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_845 <= 32'h34d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_845 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_846 <= 32'h34e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_846 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_847 <= 32'h34f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h34f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_847 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_848 <= 32'h350; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h350 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_848 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_849 <= 32'h351; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h351 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_849 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_850 <= 32'h352; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h352 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_850 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_851 <= 32'h353; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h353 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_851 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_852 <= 32'h354; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h354 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_852 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_853 <= 32'h355; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h355 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_853 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_854 <= 32'h356; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h356 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_854 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_855 <= 32'h357; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h357 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_855 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_856 <= 32'h358; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h358 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_856 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_857 <= 32'h359; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h359 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_857 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_858 <= 32'h35a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_858 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_859 <= 32'h35b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_859 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_860 <= 32'h35c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_860 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_861 <= 32'h35d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_861 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_862 <= 32'h35e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_862 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_863 <= 32'h35f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h35f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_863 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_864 <= 32'h360; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h360 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_864 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_865 <= 32'h361; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h361 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_865 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_866 <= 32'h362; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h362 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_866 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_867 <= 32'h363; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h363 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_867 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_868 <= 32'h364; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h364 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_868 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_869 <= 32'h365; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h365 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_869 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_870 <= 32'h366; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h366 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_870 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_871 <= 32'h367; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h367 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_871 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_872 <= 32'h368; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h368 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_872 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_873 <= 32'h369; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h369 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_873 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_874 <= 32'h36a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_874 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_875 <= 32'h36b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_875 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_876 <= 32'h36c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_876 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_877 <= 32'h36d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_877 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_878 <= 32'h36e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_878 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_879 <= 32'h36f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h36f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_879 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_880 <= 32'h370; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h370 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_880 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_881 <= 32'h371; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h371 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_881 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_882 <= 32'h372; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h372 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_882 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_883 <= 32'h373; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h373 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_883 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_884 <= 32'h374; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h374 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_884 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_885 <= 32'h375; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h375 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_885 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_886 <= 32'h376; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h376 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_886 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_887 <= 32'h377; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h377 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_887 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_888 <= 32'h378; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h378 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_888 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_889 <= 32'h379; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h379 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_889 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_890 <= 32'h37a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_890 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_891 <= 32'h37b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_891 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_892 <= 32'h37c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_892 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_893 <= 32'h37d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_893 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_894 <= 32'h37e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_894 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_895 <= 32'h37f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h37f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_895 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_896 <= 32'h380; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h380 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_896 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_897 <= 32'h381; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h381 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_897 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_898 <= 32'h382; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h382 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_898 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_899 <= 32'h383; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h383 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_899 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_900 <= 32'h384; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h384 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_900 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_901 <= 32'h385; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h385 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_901 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_902 <= 32'h386; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h386 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_902 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_903 <= 32'h387; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h387 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_903 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_904 <= 32'h388; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h388 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_904 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_905 <= 32'h389; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h389 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_905 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_906 <= 32'h38a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_906 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_907 <= 32'h38b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_907 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_908 <= 32'h38c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_908 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_909 <= 32'h38d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_909 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_910 <= 32'h38e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_910 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_911 <= 32'h38f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h38f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_911 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_912 <= 32'h390; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h390 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_912 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_913 <= 32'h391; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h391 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_913 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_914 <= 32'h392; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h392 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_914 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_915 <= 32'h393; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h393 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_915 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_916 <= 32'h394; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h394 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_916 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_917 <= 32'h395; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h395 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_917 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_918 <= 32'h396; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h396 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_918 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_919 <= 32'h397; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h397 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_919 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_920 <= 32'h398; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h398 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_920 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_921 <= 32'h399; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h399 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_921 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_922 <= 32'h39a; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39a == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_922 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_923 <= 32'h39b; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39b == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_923 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_924 <= 32'h39c; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39c == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_924 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_925 <= 32'h39d; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39d == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_925 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_926 <= 32'h39e; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39e == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_926 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_927 <= 32'h39f; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h39f == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_927 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_928 <= 32'h3a0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_928 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_929 <= 32'h3a1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_929 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_930 <= 32'h3a2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_930 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_931 <= 32'h3a3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_931 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_932 <= 32'h3a4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_932 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_933 <= 32'h3a5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_933 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_934 <= 32'h3a6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_934 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_935 <= 32'h3a7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_935 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_936 <= 32'h3a8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_936 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_937 <= 32'h3a9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3a9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_937 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_938 <= 32'h3aa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3aa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_938 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_939 <= 32'h3ab; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ab == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_939 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_940 <= 32'h3ac; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ac == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_940 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_941 <= 32'h3ad; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ad == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_941 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_942 <= 32'h3ae; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ae == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_942 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_943 <= 32'h3af; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3af == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_943 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_944 <= 32'h3b0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_944 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_945 <= 32'h3b1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_945 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_946 <= 32'h3b2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_946 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_947 <= 32'h3b3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_947 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_948 <= 32'h3b4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_948 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_949 <= 32'h3b5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_949 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_950 <= 32'h3b6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_950 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_951 <= 32'h3b7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_951 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_952 <= 32'h3b8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_952 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_953 <= 32'h3b9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3b9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_953 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_954 <= 32'h3ba; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ba == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_954 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_955 <= 32'h3bb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3bb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_955 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_956 <= 32'h3bc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3bc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_956 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_957 <= 32'h3bd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3bd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_957 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_958 <= 32'h3be; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3be == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_958 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_959 <= 32'h3bf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3bf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_959 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_960 <= 32'h3c0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_960 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_961 <= 32'h3c1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_961 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_962 <= 32'h3c2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_962 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_963 <= 32'h3c3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_963 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_964 <= 32'h3c4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_964 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_965 <= 32'h3c5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_965 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_966 <= 32'h3c6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_966 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_967 <= 32'h3c7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_967 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_968 <= 32'h3c8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_968 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_969 <= 32'h3c9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3c9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_969 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_970 <= 32'h3ca; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ca == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_970 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_971 <= 32'h3cb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3cb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_971 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_972 <= 32'h3cc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3cc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_972 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_973 <= 32'h3cd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3cd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_973 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_974 <= 32'h3ce; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ce == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_974 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_975 <= 32'h3cf; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3cf == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_975 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_976 <= 32'h3d0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_976 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_977 <= 32'h3d1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_977 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_978 <= 32'h3d2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_978 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_979 <= 32'h3d3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_979 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_980 <= 32'h3d4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_980 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_981 <= 32'h3d5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_981 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_982 <= 32'h3d6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_982 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_983 <= 32'h3d7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_983 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_984 <= 32'h3d8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_984 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_985 <= 32'h3d9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3d9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_985 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_986 <= 32'h3da; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3da == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_986 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_987 <= 32'h3db; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3db == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_987 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_988 <= 32'h3dc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3dc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_988 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_989 <= 32'h3dd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3dd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_989 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_990 <= 32'h3de; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3de == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_990 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_991 <= 32'h3df; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3df == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_991 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_992 <= 32'h3e0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_992 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_993 <= 32'h3e1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_993 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_994 <= 32'h3e2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_994 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_995 <= 32'h3e3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_995 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_996 <= 32'h3e4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_996 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_997 <= 32'h3e5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_997 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_998 <= 32'h3e6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_998 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_999 <= 32'h3e7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_999 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1000 <= 32'h3e8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1000 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1001 <= 32'h3e9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3e9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1001 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1002 <= 32'h3ea; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ea == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1002 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1003 <= 32'h3eb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3eb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1003 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1004 <= 32'h3ec; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ec == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1004 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1005 <= 32'h3ed; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ed == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1005 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1006 <= 32'h3ee; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ee == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1006 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1007 <= 32'h3ef; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ef == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1007 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1008 <= 32'h3f0; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f0 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1008 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1009 <= 32'h3f1; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f1 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1009 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1010 <= 32'h3f2; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f2 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1010 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1011 <= 32'h3f3; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f3 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1011 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1012 <= 32'h3f4; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f4 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1012 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1013 <= 32'h3f5; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f5 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1013 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1014 <= 32'h3f6; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f6 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1014 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1015 <= 32'h3f7; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f7 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1015 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1016 <= 32'h3f8; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f8 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1016 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1017 <= 32'h3f9; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3f9 == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1017 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1018 <= 32'h3fa; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3fa == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1018 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1019 <= 32'h3fb; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3fb == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1019 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1020 <= 32'h3fc; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3fc == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1020 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1021 <= 32'h3fd; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3fd == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1021 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1022 <= 32'h3fe; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3fe == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1022 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (reset) begin // @[DataMemoryTest.scala 16:20]
      mem_1023 <= 32'h3ff; // @[DataMemoryTest.scala 16:20]
    end else if (io_enableWrite) begin // @[DataMemoryTest.scala 22:23]
      if (10'h3ff == io_addr) begin // @[DataMemoryTest.scala 23:18]
        mem_1023 <= io_dataIn; // @[DataMemoryTest.scala 23:18]
      end
    end
    if (10'h3ff == io_addr) begin // @[DataMemoryTest.scala 19:24]
      io_dataOut_REG <= mem_1023; // @[DataMemoryTest.scala 19:24]
    end else if (10'h3fe == io_addr) begin // @[DataMemoryTest.scala 19:24]
      io_dataOut_REG <= mem_1022; // @[DataMemoryTest.scala 19:24]
    end else if (10'h3fd == io_addr) begin // @[DataMemoryTest.scala 19:24]
      io_dataOut_REG <= mem_1021; // @[DataMemoryTest.scala 19:24]
    end else if (10'h3fc == io_addr) begin // @[DataMemoryTest.scala 19:24]
      io_dataOut_REG <= mem_1020; // @[DataMemoryTest.scala 19:24]
    end else begin
      io_dataOut_REG <= _GEN_1019;
    end
    io_dataOut_REG_1 <= io_dataIn; // @[DataMemoryTest.scala 24:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mem_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mem_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mem_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mem_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mem_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mem_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mem_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mem_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mem_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mem_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mem_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mem_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mem_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mem_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mem_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mem_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mem_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mem_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mem_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mem_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mem_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mem_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mem_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mem_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mem_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mem_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mem_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  mem_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  mem_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  mem_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  mem_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  mem_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  mem_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  mem_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  mem_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  mem_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  mem_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  mem_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  mem_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  mem_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  mem_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  mem_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  mem_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  mem_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  mem_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  mem_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  mem_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  mem_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  mem_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  mem_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  mem_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  mem_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  mem_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  mem_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  mem_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  mem_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  mem_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  mem_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  mem_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  mem_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  mem_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  mem_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  mem_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  mem_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  mem_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  mem_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  mem_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  mem_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  mem_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  mem_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  mem_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  mem_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  mem_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  mem_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  mem_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  mem_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  mem_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  mem_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  mem_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  mem_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  mem_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  mem_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  mem_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  mem_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  mem_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  mem_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  mem_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  mem_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  mem_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  mem_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  mem_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  mem_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  mem_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  mem_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  mem_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  mem_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  mem_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  mem_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  mem_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  mem_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  mem_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  mem_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  mem_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  mem_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  mem_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  mem_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  mem_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  mem_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  mem_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  mem_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  mem_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  mem_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  mem_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  mem_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  mem_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  mem_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  mem_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  mem_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  mem_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  mem_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  mem_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  mem_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  mem_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  mem_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  mem_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  mem_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  mem_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  mem_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  mem_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  mem_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  mem_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  mem_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  mem_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  mem_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  mem_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  mem_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  mem_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  mem_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  mem_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  mem_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  mem_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  mem_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  mem_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  mem_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  mem_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  mem_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  mem_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  mem_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  mem_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  mem_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  mem_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  mem_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  mem_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  mem_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  mem_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  mem_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  mem_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  mem_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  mem_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  mem_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  mem_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  mem_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  mem_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  mem_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  mem_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  mem_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  mem_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  mem_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  mem_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  mem_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  mem_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  mem_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  mem_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  mem_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  mem_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  mem_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  mem_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  mem_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  mem_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  mem_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  mem_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  mem_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  mem_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  mem_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  mem_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  mem_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  mem_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  mem_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  mem_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  mem_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  mem_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  mem_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  mem_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  mem_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  mem_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  mem_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  mem_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  mem_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  mem_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  mem_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  mem_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  mem_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  mem_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  mem_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  mem_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  mem_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  mem_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  mem_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  mem_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  mem_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  mem_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  mem_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  mem_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  mem_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  mem_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  mem_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  mem_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  mem_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  mem_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  mem_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  mem_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  mem_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  mem_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  mem_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  mem_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  mem_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  mem_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  mem_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  mem_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  mem_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  mem_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  mem_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  mem_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  mem_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  mem_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  mem_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  mem_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  mem_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  mem_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  mem_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  mem_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  mem_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  mem_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  mem_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  mem_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  mem_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  mem_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  mem_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  mem_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  mem_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  mem_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  mem_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  mem_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  mem_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  mem_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  mem_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  mem_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  mem_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  mem_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  mem_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  mem_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  mem_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  mem_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  mem_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  mem_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  mem_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  mem_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  mem_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  mem_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  mem_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  mem_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  mem_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  mem_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  mem_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  mem_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  mem_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  mem_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  mem_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  mem_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  mem_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  mem_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  mem_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  mem_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  mem_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  mem_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  mem_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  mem_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  mem_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  mem_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  mem_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  mem_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  mem_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  mem_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  mem_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  mem_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  mem_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  mem_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  mem_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  mem_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  mem_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  mem_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  mem_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  mem_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  mem_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  mem_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  mem_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  mem_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  mem_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  mem_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  mem_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  mem_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  mem_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  mem_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  mem_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  mem_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  mem_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  mem_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  mem_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  mem_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  mem_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  mem_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  mem_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  mem_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  mem_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  mem_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  mem_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  mem_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  mem_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  mem_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  mem_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  mem_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  mem_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  mem_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  mem_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  mem_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  mem_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  mem_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  mem_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  mem_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  mem_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  mem_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  mem_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  mem_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  mem_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  mem_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  mem_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  mem_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  mem_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  mem_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  mem_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  mem_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  mem_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  mem_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  mem_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  mem_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  mem_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  mem_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  mem_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  mem_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  mem_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  mem_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  mem_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  mem_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  mem_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  mem_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  mem_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  mem_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  mem_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  mem_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  mem_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  mem_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  mem_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  mem_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  mem_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  mem_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  mem_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  mem_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  mem_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  mem_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  mem_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  mem_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  mem_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  mem_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  mem_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  mem_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  mem_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  mem_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  mem_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  mem_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  mem_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  mem_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  mem_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  mem_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  mem_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  mem_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  mem_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  mem_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  mem_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  mem_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  mem_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  mem_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  mem_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  mem_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  mem_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  mem_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  mem_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  mem_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  mem_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  mem_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  mem_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  mem_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  mem_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  mem_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  mem_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  mem_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  mem_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  mem_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  mem_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  mem_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  mem_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  mem_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  mem_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  mem_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  mem_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  mem_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  mem_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  mem_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  mem_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  mem_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  mem_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  mem_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  mem_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  mem_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  mem_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  mem_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  mem_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  mem_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  mem_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  mem_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  mem_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  mem_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  mem_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  mem_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  mem_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  mem_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  mem_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  mem_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  mem_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  mem_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  mem_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  mem_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  mem_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  mem_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  mem_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  mem_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  mem_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  mem_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  mem_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  mem_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  mem_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  mem_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  mem_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  mem_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  mem_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  mem_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  mem_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  mem_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  mem_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  mem_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  mem_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  mem_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  mem_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  mem_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  mem_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  mem_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  mem_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  mem_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  mem_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  mem_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  mem_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  mem_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  mem_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  mem_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  mem_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  mem_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  mem_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  mem_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  mem_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  mem_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  mem_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  mem_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  mem_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  mem_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  mem_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  mem_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  mem_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  mem_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  mem_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  mem_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  mem_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  mem_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  mem_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  mem_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  mem_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  mem_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  mem_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  mem_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  mem_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  mem_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  mem_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  mem_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  mem_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  mem_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  mem_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  mem_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  mem_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  mem_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  mem_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  mem_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  mem_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  mem_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  mem_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  mem_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  mem_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  mem_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  mem_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  mem_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  mem_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  mem_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  mem_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  mem_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  mem_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  mem_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  mem_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  mem_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  mem_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  mem_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  mem_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  mem_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  mem_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  mem_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  mem_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  mem_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  mem_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  mem_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  mem_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  mem_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  mem_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  mem_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  mem_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  mem_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  mem_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  mem_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  mem_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  mem_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  mem_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  mem_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  mem_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  mem_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  mem_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  mem_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  mem_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  mem_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  mem_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  mem_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  mem_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  mem_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  mem_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  mem_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  mem_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  mem_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  mem_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  mem_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  mem_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  mem_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  mem_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  mem_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  mem_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  mem_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  mem_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  mem_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  mem_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  mem_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  mem_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  mem_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  mem_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  mem_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  mem_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  mem_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  mem_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  mem_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  mem_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  mem_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  mem_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  mem_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  mem_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  mem_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  mem_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  mem_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  mem_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  mem_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  mem_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  mem_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  mem_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  mem_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  mem_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  mem_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  mem_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  mem_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  mem_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  mem_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  mem_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  mem_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  mem_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  mem_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  mem_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  mem_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  mem_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  mem_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  mem_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  mem_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  mem_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  mem_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  mem_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  mem_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  mem_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  mem_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  mem_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  mem_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  mem_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  mem_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  mem_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  mem_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  mem_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  mem_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  mem_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  mem_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  mem_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  mem_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  mem_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  mem_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  mem_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  mem_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  mem_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  mem_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  mem_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  mem_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  mem_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  mem_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  mem_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  mem_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  mem_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  mem_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  mem_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  mem_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  mem_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  mem_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  mem_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  mem_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  mem_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  mem_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  mem_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  mem_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  mem_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  mem_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  mem_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  mem_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  mem_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  mem_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  mem_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  mem_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  mem_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  mem_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  mem_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  mem_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  mem_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  mem_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  mem_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  mem_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  mem_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  mem_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  mem_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  mem_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  mem_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  mem_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  mem_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  mem_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  mem_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  mem_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  mem_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  mem_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  mem_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  mem_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  mem_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  mem_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  mem_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  mem_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  mem_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  mem_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  mem_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  mem_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  mem_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  mem_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  mem_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  mem_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  mem_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  mem_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  mem_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  mem_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  mem_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  mem_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  mem_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  mem_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  mem_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  mem_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  mem_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  mem_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  mem_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  mem_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  mem_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  mem_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  mem_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  mem_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  mem_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  mem_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  mem_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  mem_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  mem_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  mem_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  mem_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  mem_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  mem_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  mem_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  mem_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  mem_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  mem_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  mem_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  mem_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  mem_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  mem_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  mem_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  mem_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  mem_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  mem_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  mem_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  mem_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  mem_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  mem_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  mem_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  mem_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  mem_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  mem_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  mem_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  mem_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  mem_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  mem_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  mem_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  mem_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  mem_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  mem_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  mem_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  mem_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  mem_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  mem_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  mem_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  mem_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  mem_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  mem_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  mem_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  mem_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  mem_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  mem_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  mem_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  mem_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  mem_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  mem_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  mem_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  mem_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  mem_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  mem_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  mem_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  mem_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  mem_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  mem_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  mem_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  mem_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  mem_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  mem_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  mem_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  mem_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  mem_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  mem_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  mem_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  mem_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  mem_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  mem_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  mem_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  mem_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  mem_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  mem_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  mem_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  mem_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  mem_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  mem_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  mem_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  mem_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  mem_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  mem_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  mem_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  mem_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  mem_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  mem_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  mem_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  mem_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  mem_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  mem_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  mem_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  mem_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  mem_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  mem_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  mem_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  mem_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  mem_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  mem_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  mem_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  mem_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  mem_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  mem_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  mem_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  mem_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  mem_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  mem_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  mem_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  mem_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  mem_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  mem_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  mem_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  mem_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  mem_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  mem_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  mem_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  mem_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  mem_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  mem_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  mem_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  mem_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  mem_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  mem_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  mem_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  mem_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  mem_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  mem_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  mem_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  mem_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  mem_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  mem_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  mem_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  mem_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  mem_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  mem_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  mem_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  mem_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  mem_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  mem_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  mem_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  mem_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  mem_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  mem_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  mem_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  mem_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  mem_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  mem_999 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  mem_1000 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  mem_1001 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  mem_1002 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  mem_1003 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  mem_1004 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  mem_1005 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  mem_1006 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  mem_1007 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  mem_1008 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  mem_1009 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  mem_1010 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  mem_1011 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  mem_1012 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  mem_1013 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  mem_1014 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  mem_1015 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  mem_1016 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  mem_1017 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  mem_1018 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  mem_1019 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  mem_1020 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  mem_1021 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  mem_1022 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  mem_1023 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  io_dataOut_REG = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  io_dataOut_REG_1 = _RAND_1025[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemoryMappedLeds(
  input         clock,
  input         reset,
  input         io_port_write,
  input  [31:0] io_port_wrData,
  output [31:0] io_port_rdData,
  output [15:0] io_pins
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ledReg; // @[MemoryMappedLeds.scala 28:23]
  wire [31:0] _GEN_0 = io_port_write ? io_port_wrData : {{16'd0}, ledReg}; // @[MemoryMappedLeds.scala 30:23 31:12 28:23]
  wire [31:0] _GEN_1 = reset ? 32'h0 : _GEN_0; // @[MemoryMappedLeds.scala 28:{23,23}]
  assign io_port_rdData = {{16'd0}, ledReg}; // @[MemoryMappedLeds.scala 35:18]
  assign io_pins = ledReg; // @[MemoryMappedLeds.scala 34:11]
  always @(posedge clock) begin
    ledReg <= _GEN_1[15:0]; // @[MemoryMappedLeds.scala 28:{23,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ledReg = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemoryMappedIO(
  input         clock,
  input         reset,
  input  [31:0] io_address,
  input  [31:0] io_dataWriteMem,
  input         io_writeEnable,
  output [31:0] io_dataReadIO,
  output [15:0] io_leds
);
  wire  leds_clock; // @[MemoryMappedIO.scala 21:20]
  wire  leds_reset; // @[MemoryMappedIO.scala 21:20]
  wire  leds_io_port_write; // @[MemoryMappedIO.scala 21:20]
  wire [31:0] leds_io_port_wrData; // @[MemoryMappedIO.scala 21:20]
  wire [31:0] leds_io_port_rdData; // @[MemoryMappedIO.scala 21:20]
  wire [15:0] leds_io_pins; // @[MemoryMappedIO.scala 21:20]
  wire [31:0] addressIO = io_address - 32'h400; // @[MemoryMappedIO.scala 24:30]
  MemoryMappedLeds leds ( // @[MemoryMappedIO.scala 21:20]
    .clock(leds_clock),
    .reset(leds_reset),
    .io_port_write(leds_io_port_write),
    .io_port_wrData(leds_io_port_wrData),
    .io_port_rdData(leds_io_port_rdData),
    .io_pins(leds_io_pins)
  );
  assign io_dataReadIO = leds_io_port_rdData; // @[MemoryMappedIO.scala 32:17]
  assign io_leds = leds_io_pins; // @[MemoryMappedIO.scala 33:11]
  assign leds_clock = clock;
  assign leds_reset = reset;
  assign leds_io_port_write = io_writeEnable & addressIO == 32'h0; // @[MemoryMappedIO.scala 28:40]
  assign leds_io_port_wrData = {{16'd0}, io_dataWriteMem[15:0]}; // @[MemoryMappedIO.scala 29:23]
endmodule
module MEMStage(
  input         clock,
  input         reset,
  input  [31:0] io_ALURes,
  input  [31:0] io_address,
  input  [31:0] io_dataWriteMem,
  input         io_memWriteEnable,
  input         io_registerWriteEnableIn,
  input         io_writeDataMux,
  input  [4:0]  io_rdRegIn,
  input         io_readIsIO,
  input         io_IOWriteEnable,
  output [31:0] io_writeData,
  output        io_registerWriteEnableOut,
  output [4:0]  io_rdRegOut,
  output [15:0] io_leds
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  dataMem_clock; // @[MEMStage.scala 36:23]
  wire  dataMem_reset; // @[MEMStage.scala 36:23]
  wire [9:0] dataMem_io_addr; // @[MEMStage.scala 36:23]
  wire  dataMem_io_enableWrite; // @[MEMStage.scala 36:23]
  wire [31:0] dataMem_io_dataIn; // @[MEMStage.scala 36:23]
  wire [31:0] dataMem_io_dataOut; // @[MEMStage.scala 36:23]
  wire  memoryMappedIO_clock; // @[MEMStage.scala 41:30]
  wire  memoryMappedIO_reset; // @[MEMStage.scala 41:30]
  wire [31:0] memoryMappedIO_io_address; // @[MEMStage.scala 41:30]
  wire [31:0] memoryMappedIO_io_dataWriteMem; // @[MEMStage.scala 41:30]
  wire  memoryMappedIO_io_writeEnable; // @[MEMStage.scala 41:30]
  wire [31:0] memoryMappedIO_io_dataReadIO; // @[MEMStage.scala 41:30]
  wire [15:0] memoryMappedIO_io_leds; // @[MEMStage.scala 41:30]
  reg [31:0] ALUResReg; // @[MEMStage.scala 33:26]
  reg [1:0] controlReg; // @[MEMStage.scala 34:27]
  reg [4:0] rdReg; // @[MEMStage.scala 35:22]
  reg  readIsIO; // @[MEMStage.scala 38:25]
  wire [1:0] _controlReg_T = {io_registerWriteEnableIn,io_writeDataMux}; // @[Cat.scala 33:92]
  wire [31:0] _io_writeData_T = readIsIO ? memoryMappedIO_io_dataReadIO : dataMem_io_dataOut; // @[MEMStage.scala 55:24]
  DataMemoryTest dataMem ( // @[MEMStage.scala 36:23]
    .clock(dataMem_clock),
    .reset(dataMem_reset),
    .io_addr(dataMem_io_addr),
    .io_enableWrite(dataMem_io_enableWrite),
    .io_dataIn(dataMem_io_dataIn),
    .io_dataOut(dataMem_io_dataOut)
  );
  MemoryMappedIO memoryMappedIO ( // @[MEMStage.scala 41:30]
    .clock(memoryMappedIO_clock),
    .reset(memoryMappedIO_reset),
    .io_address(memoryMappedIO_io_address),
    .io_dataWriteMem(memoryMappedIO_io_dataWriteMem),
    .io_writeEnable(memoryMappedIO_io_writeEnable),
    .io_dataReadIO(memoryMappedIO_io_dataReadIO),
    .io_leds(memoryMappedIO_io_leds)
  );
  assign io_writeData = controlReg[0] ? _io_writeData_T : ALUResReg; // @[MEMStage.scala 54:30 55:18 57:18]
  assign io_registerWriteEnableOut = controlReg[1]; // @[MEMStage.scala 59:42]
  assign io_rdRegOut = rdReg; // @[MEMStage.scala 60:15]
  assign io_leds = memoryMappedIO_io_leds; // @[MEMStage.scala 45:11]
  assign dataMem_clock = clock;
  assign dataMem_reset = reset;
  assign dataMem_io_addr = io_address[9:0]; // @[MEMStage.scala 64:19]
  assign dataMem_io_enableWrite = io_memWriteEnable; // @[MEMStage.scala 66:26]
  assign dataMem_io_dataIn = io_dataWriteMem; // @[MEMStage.scala 65:21]
  assign memoryMappedIO_clock = clock;
  assign memoryMappedIO_reset = reset;
  assign memoryMappedIO_io_address = io_address; // @[MEMStage.scala 44:29]
  assign memoryMappedIO_io_dataWriteMem = io_dataWriteMem; // @[MEMStage.scala 43:34]
  assign memoryMappedIO_io_writeEnable = io_IOWriteEnable; // @[MEMStage.scala 42:33]
  always @(posedge clock) begin
    if (reset) begin // @[MEMStage.scala 33:26]
      ALUResReg <= 32'h0; // @[MEMStage.scala 33:26]
    end else begin
      ALUResReg <= io_ALURes; // @[MEMStage.scala 48:13]
    end
    if (reset) begin // @[MEMStage.scala 34:27]
      controlReg <= 2'h0; // @[MEMStage.scala 34:27]
    end else begin
      controlReg <= _controlReg_T; // @[MEMStage.scala 49:14]
    end
    if (reset) begin // @[MEMStage.scala 35:22]
      rdReg <= 5'h0; // @[MEMStage.scala 35:22]
    end else begin
      rdReg <= io_rdRegIn; // @[MEMStage.scala 50:9]
    end
    readIsIO <= io_readIsIO; // @[MEMStage.scala 38:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ALUResReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  controlReg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rdReg = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  readIsIO = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ProcessorTopLevel(
  input         clock,
  input         reset,
  output [15:0] io_LEDs
);
  wire  IF_clock; // @[ProcessorTopLevel.scala 14:18]
  wire  IF_reset; // @[ProcessorTopLevel.scala 14:18]
  wire [31:0] IF_io_instruction; // @[ProcessorTopLevel.scala 14:18]
  wire [31:0] ID_io_instruction; // @[ProcessorTopLevel.scala 15:18]
  wire [4:0] ID_io_rs1; // @[ProcessorTopLevel.scala 15:18]
  wire [4:0] ID_io_rs2; // @[ProcessorTopLevel.scala 15:18]
  wire [4:0] ID_io_rd; // @[ProcessorTopLevel.scala 15:18]
  wire [2:0] ID_io_funct3; // @[ProcessorTopLevel.scala 15:18]
  wire [6:0] ID_io_funct7; // @[ProcessorTopLevel.scala 15:18]
  wire [2:0] ID_io_instrType; // @[ProcessorTopLevel.scala 15:18]
  wire [6:0] ID_io_opcode; // @[ProcessorTopLevel.scala 15:18]
  wire  EX_clock; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_reset; // @[ProcessorTopLevel.scala 16:18]
  wire [31:0] EX_io_instruction; // @[ProcessorTopLevel.scala 16:18]
  wire [2:0] EX_io_instrType; // @[ProcessorTopLevel.scala 16:18]
  wire [2:0] EX_io_funct3; // @[ProcessorTopLevel.scala 16:18]
  wire [6:0] EX_io_funct7; // @[ProcessorTopLevel.scala 16:18]
  wire [6:0] EX_io_opcode; // @[ProcessorTopLevel.scala 16:18]
  wire [4:0] EX_io_rs1; // @[ProcessorTopLevel.scala 16:18]
  wire [4:0] EX_io_rs2; // @[ProcessorTopLevel.scala 16:18]
  wire [4:0] EX_io_rd; // @[ProcessorTopLevel.scala 16:18]
  wire [31:0] EX_io_writeData; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_writeEnable; // @[ProcessorTopLevel.scala 16:18]
  wire [4:0] EX_io_rdReg; // @[ProcessorTopLevel.scala 16:18]
  wire [31:0] EX_io_ALURes; // @[ProcessorTopLevel.scala 16:18]
  wire [31:0] EX_io_address; // @[ProcessorTopLevel.scala 16:18]
  wire [31:0] EX_io_dataWriteMem; // @[ProcessorTopLevel.scala 16:18]
  wire [4:0] EX_io_rdRegIn; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_RegWriteEnable; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_WriteDataMux; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_MemWriteEnable; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_readIsIO; // @[ProcessorTopLevel.scala 16:18]
  wire  EX_io_IOWriteEnable; // @[ProcessorTopLevel.scala 16:18]
  wire  MEM_clock; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_reset; // @[ProcessorTopLevel.scala 17:20]
  wire [31:0] MEM_io_ALURes; // @[ProcessorTopLevel.scala 17:20]
  wire [31:0] MEM_io_address; // @[ProcessorTopLevel.scala 17:20]
  wire [31:0] MEM_io_dataWriteMem; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_memWriteEnable; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_registerWriteEnableIn; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_writeDataMux; // @[ProcessorTopLevel.scala 17:20]
  wire [4:0] MEM_io_rdRegIn; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_readIsIO; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_IOWriteEnable; // @[ProcessorTopLevel.scala 17:20]
  wire [31:0] MEM_io_writeData; // @[ProcessorTopLevel.scala 17:20]
  wire  MEM_io_registerWriteEnableOut; // @[ProcessorTopLevel.scala 17:20]
  wire [4:0] MEM_io_rdRegOut; // @[ProcessorTopLevel.scala 17:20]
  wire [15:0] MEM_io_leds; // @[ProcessorTopLevel.scala 17:20]
  IFStage IF ( // @[ProcessorTopLevel.scala 14:18]
    .clock(IF_clock),
    .reset(IF_reset),
    .io_instruction(IF_io_instruction)
  );
  InstructionDecoder ID ( // @[ProcessorTopLevel.scala 15:18]
    .io_instruction(ID_io_instruction),
    .io_rs1(ID_io_rs1),
    .io_rs2(ID_io_rs2),
    .io_rd(ID_io_rd),
    .io_funct3(ID_io_funct3),
    .io_funct7(ID_io_funct7),
    .io_instrType(ID_io_instrType),
    .io_opcode(ID_io_opcode)
  );
  EXStage EX ( // @[ProcessorTopLevel.scala 16:18]
    .clock(EX_clock),
    .reset(EX_reset),
    .io_instruction(EX_io_instruction),
    .io_instrType(EX_io_instrType),
    .io_funct3(EX_io_funct3),
    .io_funct7(EX_io_funct7),
    .io_opcode(EX_io_opcode),
    .io_rs1(EX_io_rs1),
    .io_rs2(EX_io_rs2),
    .io_rd(EX_io_rd),
    .io_writeData(EX_io_writeData),
    .io_writeEnable(EX_io_writeEnable),
    .io_rdReg(EX_io_rdReg),
    .io_ALURes(EX_io_ALURes),
    .io_address(EX_io_address),
    .io_dataWriteMem(EX_io_dataWriteMem),
    .io_rdRegIn(EX_io_rdRegIn),
    .io_RegWriteEnable(EX_io_RegWriteEnable),
    .io_WriteDataMux(EX_io_WriteDataMux),
    .io_MemWriteEnable(EX_io_MemWriteEnable),
    .io_readIsIO(EX_io_readIsIO),
    .io_IOWriteEnable(EX_io_IOWriteEnable)
  );
  MEMStage MEM ( // @[ProcessorTopLevel.scala 17:20]
    .clock(MEM_clock),
    .reset(MEM_reset),
    .io_ALURes(MEM_io_ALURes),
    .io_address(MEM_io_address),
    .io_dataWriteMem(MEM_io_dataWriteMem),
    .io_memWriteEnable(MEM_io_memWriteEnable),
    .io_registerWriteEnableIn(MEM_io_registerWriteEnableIn),
    .io_writeDataMux(MEM_io_writeDataMux),
    .io_rdRegIn(MEM_io_rdRegIn),
    .io_readIsIO(MEM_io_readIsIO),
    .io_IOWriteEnable(MEM_io_IOWriteEnable),
    .io_writeData(MEM_io_writeData),
    .io_registerWriteEnableOut(MEM_io_registerWriteEnableOut),
    .io_rdRegOut(MEM_io_rdRegOut),
    .io_leds(MEM_io_leds)
  );
  assign io_LEDs = MEM_io_leds; // @[ProcessorTopLevel.scala 54:11]
  assign IF_clock = clock;
  assign IF_reset = reset;
  assign ID_io_instruction = IF_io_instruction; // @[ProcessorTopLevel.scala 22:21]
  assign EX_clock = clock;
  assign EX_reset = reset;
  assign EX_io_instruction = IF_io_instruction; // @[ProcessorTopLevel.scala 25:21]
  assign EX_io_instrType = ID_io_instrType; // @[ProcessorTopLevel.scala 26:19]
  assign EX_io_funct3 = ID_io_funct3; // @[ProcessorTopLevel.scala 27:16]
  assign EX_io_funct7 = ID_io_funct7; // @[ProcessorTopLevel.scala 28:16]
  assign EX_io_opcode = ID_io_opcode; // @[ProcessorTopLevel.scala 29:16]
  assign EX_io_rs1 = ID_io_rs1; // @[ProcessorTopLevel.scala 30:13]
  assign EX_io_rs2 = ID_io_rs2; // @[ProcessorTopLevel.scala 31:13]
  assign EX_io_rd = ID_io_rd; // @[ProcessorTopLevel.scala 32:12]
  assign EX_io_writeData = MEM_io_writeData; // @[ProcessorTopLevel.scala 46:19]
  assign EX_io_writeEnable = MEM_io_registerWriteEnableOut; // @[ProcessorTopLevel.scala 47:21]
  assign EX_io_rdReg = MEM_io_rdRegOut; // @[ProcessorTopLevel.scala 48:15]
  assign MEM_clock = clock;
  assign MEM_reset = reset;
  assign MEM_io_ALURes = EX_io_ALURes; // @[ProcessorTopLevel.scala 35:17]
  assign MEM_io_address = EX_io_address; // @[ProcessorTopLevel.scala 36:18]
  assign MEM_io_dataWriteMem = EX_io_dataWriteMem; // @[ProcessorTopLevel.scala 37:23]
  assign MEM_io_memWriteEnable = EX_io_MemWriteEnable; // @[ProcessorTopLevel.scala 38:25]
  assign MEM_io_registerWriteEnableIn = EX_io_RegWriteEnable; // @[ProcessorTopLevel.scala 39:32]
  assign MEM_io_writeDataMux = EX_io_WriteDataMux; // @[ProcessorTopLevel.scala 40:23]
  assign MEM_io_rdRegIn = EX_io_rdRegIn; // @[ProcessorTopLevel.scala 41:18]
  assign MEM_io_readIsIO = EX_io_readIsIO; // @[ProcessorTopLevel.scala 44:19]
  assign MEM_io_IOWriteEnable = EX_io_IOWriteEnable; // @[ProcessorTopLevel.scala 43:24]
endmodule
